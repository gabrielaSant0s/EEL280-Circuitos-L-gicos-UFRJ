CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 949 95 0 1 11
0 19
0
0 0 21360 270
2 0V
-7 -23 7 -15
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6369 0 0
2
5.89916e-315 0
0
5 4073~
219 167 519 0 4 22
0 6 5 4 3
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 9 0
1 U
9172 0 0
2
43788.1 0
0
6 74LS48
188 311 678 0 14 29
0 2 9 8 7 33 34 16 15 14
13 12 11 10 35
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
3 U13
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7100 0 0
2
43788.1 0
0
7 Ground~
168 243 600 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
43788.1 1
0
9 CC 7-Seg~
183 434 585 0 17 19
10 10 11 12 13 14 15 16 36 2
0 0 1 1 1 1 1 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7678 0 0
2
43788.1 2
0
7 Ground~
168 434 528 0 1 3
0 2
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
961 0 0
2
43788.1 3
0
5 4082~
219 750 620 0 5 22
0 18 19 5 20 21
0
0 0 624 180
4 4082
-7 -24 21 -16
3 U5A
-13 -28 8 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
3178 0 0
2
43788.1 4
0
5 4071~
219 681 720 0 3 22
0 24 25 7
0
0 0 624 180
4 4071
-7 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3409 0 0
2
43788.1 5
0
5 4082~
219 746 747 0 5 22
0 18 19 22 20 24
0
0 0 624 180
4 4082
-7 -24 21 -16
3 U4B
-13 -28 8 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3951 0 0
2
43788.1 6
0
5 4082~
219 745 700 0 5 22
0 18 19 23 20 25
0
0 0 624 180
4 4082
-7 -24 21 -16
3 U4A
-13 -28 8 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
8885 0 0
2
43788.1 7
0
5 4081~
219 751 575 0 3 22
0 23 18 26
0
0 0 624 180
4 4081
-7 -24 21 -16
3 U1B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
3780 0 0
2
43788.1 8
0
5 4071~
219 686 597 0 3 22
0 21 26 8
0
0 0 624 180
4 4071
-7 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
9265 0 0
2
43788.1 9
0
5 4081~
219 747 496 0 3 22
0 22 18 9
0
0 0 624 180
4 4081
-7 -24 21 -16
3 U1A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9442 0 0
2
43788.1 10
0
2 +V
167 1014 455 0 1 3
0 20
0
0 0 53744 0
2 5V
-8 -22 6 -14
2 V1
-8 -32 6 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9424 0 0
2
43788.1 11
0
14 Logic Display~
6 669 326 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.89916e-315 5.3568e-315
0
14 Logic Display~
6 543 328 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89916e-315 5.36716e-315
0
14 Logic Display~
6 403 331 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89916e-315 5.37752e-315
0
5 4027~
219 613 431 0 7 32
0 37 30 5 30 3 18 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U7A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
7168 0 0
2
5.89916e-315 5.38788e-315
0
9 Inverter~
13 981 138 0 2 22
0 19 28
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U8A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3171 0 0
2
5.89916e-315 5.39306e-315
0
14 Logic Display~
6 193 311 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.89916e-315 5.39824e-315
0
7 Pulser~
4 153 395 0 10 12
0 38 39 40 31 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6435 0 0
2
5.89916e-315 5.40342e-315
0
5 4027~
219 344 436 0 7 32
0 41 32 31 32 3 6 23
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
5283 0 0
2
5.89916e-315 5.4086e-315
0
5 4027~
219 488 432 0 7 32
0 42 29 6 29 3 5 22
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
6874 0 0
2
5.89916e-315 5.41378e-315
0
62
0 5 3 0 0 4096 0 0 18 2 0 3
485 519
613 519
613 437
0 5 3 0 0 4096 0 0 23 3 0 3
342 519
488 519
488 438
4 5 3 0 0 4224 0 2 22 0 0 3
188 519
344 519
344 442
0 3 4 0 0 8192 0 0 2 52 0 5
650 395
650 461
84 461
84 528
143 528
0 2 5 0 0 8192 0 0 2 48 0 5
526 414
526 490
127 490
127 519
143 519
0 1 6 0 0 8192 0 0 2 50 0 5
384 418
384 474
115 474
115 510
143 510
3 4 7 0 0 8320 0 8 3 0 0 5
654 720
654 930
275 930
275 669
279 669
3 3 8 0 0 12416 0 12 3 0 0 6
659 597
581 597
581 900
260 900
260 660
279 660
3 2 9 0 0 8320 0 13 3 0 0 6
720 496
547 496
547 860
247 860
247 651
279 651
13 1 10 0 0 8320 0 3 5 0 0 3
343 696
413 696
413 621
12 2 11 0 0 4224 0 3 5 0 0 3
343 687
419 687
419 621
11 3 12 0 0 4224 0 3 5 0 0 3
343 678
425 678
425 621
10 4 13 0 0 4224 0 3 5 0 0 3
343 669
431 669
431 621
9 5 14 0 0 4224 0 3 5 0 0 3
343 660
437 660
437 621
8 6 15 0 0 4224 0 3 5 0 0 3
343 651
443 651
443 621
7 7 16 0 0 4224 0 3 5 0 0 3
343 642
449 642
449 621
1 9 2 0 0 4096 0 6 5 0 0 4
434 536
434 551
434 551
434 543
1 1 2 0 0 4224 0 3 4 0 0 3
279 642
243 642
243 608
0 0 17 0 0 8320 0 0 0 0 0 3
725 499
725 500
719 500
1 0 18 0 0 4096 0 7 0 0 46 2
768 633
902 633
2 0 19 0 0 4096 0 7 0 0 57 2
768 624
949 624
3 0 5 0 0 0 0 7 0 0 48 2
768 615
852 615
4 0 20 0 0 4096 0 7 0 0 44 2
768 606
1014 606
5 0 21 0 0 4096 0 7 0 0 38 2
723 620
721 620
1 0 18 0 0 4096 0 9 0 0 46 2
764 760
902 760
2 0 19 0 0 4096 0 9 0 0 57 2
764 751
949 751
3 0 22 0 0 4096 0 9 0 0 49 2
764 742
831 742
1 0 18 0 0 4096 0 10 0 0 46 2
763 713
902 713
2 0 19 0 0 4096 0 10 0 0 57 2
763 704
949 704
3 0 23 0 0 4096 0 10 0 0 51 2
763 695
781 695
0 2 19 0 0 0 0 0 9 0 0 3
757 752
757 751
764 751
4 0 20 0 0 4096 0 9 0 0 44 2
764 733
1014 733
4 0 20 0 0 4096 0 10 0 0 44 2
763 686
1014 686
1 5 24 0 0 8320 0 8 9 0 0 3
700 729
700 747
719 747
2 5 25 0 0 8320 0 8 10 0 0 3
700 711
700 700
718 700
1 0 23 0 0 0 0 11 0 0 51 2
769 584
781 584
2 0 18 0 0 0 0 11 0 0 46 2
769 566
902 566
1 0 21 0 0 4224 0 12 0 0 0 4
705 606
721 606
721 620
725 620
2 3 26 0 0 8320 0 12 11 0 0 3
705 588
705 575
724 575
1 0 22 0 0 0 0 13 0 0 49 2
765 505
831 505
2 0 18 0 0 0 0 13 0 0 46 2
765 487
902 487
0 3 5 0 0 0 0 0 18 48 0 2
564 404
589 404
0 3 6 0 0 0 0 0 23 50 0 3
439 406
439 405
464 405
1 0 20 0 0 4224 0 14 0 0 0 2
1014 464
1014 971
0 0 27 0 0 0 0 0 0 0 0 2
855 962
855 962
6 0 18 0 0 16512 0 18 0 0 0 5
643 413
766 413
766 196
902 196
902 976
0 0 4 0 0 16512 0 0 0 52 0 5
669 386
752 386
752 172
882 172
882 977
6 0 5 0 0 16512 0 23 0 0 0 5
518 414
564 414
564 156
852 156
852 976
1 0 22 0 0 16512 0 16 0 0 0 5
543 346
575 346
575 134
831 134
831 976
6 0 6 0 0 16512 0 22 0 0 0 5
374 418
439 418
439 121
804 121
804 972
0 0 23 0 0 16512 0 0 0 54 0 5
403 361
427 361
427 114
781 114
781 974
7 1 4 0 0 0 0 18 15 0 0 3
637 395
669 395
669 344
7 1 22 0 0 0 0 23 16 0 0 3
512 396
543 396
543 346
7 1 23 0 0 0 0 22 17 0 0 3
368 400
403 400
403 349
1 0 19 0 0 0 0 19 0 0 57 2
984 120
949 120
2 0 28 0 0 12416 0 19 0 0 0 4
984 156
984 495
985 495
985 976
1 0 19 0 0 4224 0 1 0 0 0 2
949 107
949 972
2 4 29 0 0 8320 0 23 23 0 0 4
464 396
454 396
454 414
464 414
2 4 30 0 0 12416 0 18 18 0 0 6
589 395
589 394
578 394
578 412
589 412
589 413
1 0 31 0 0 4096 0 20 0 0 61 2
193 329
193 407
3 4 31 0 0 4224 0 22 21 0 0 5
320 409
193 409
193 407
183 407
183 395
2 4 32 0 0 8320 0 22 22 0 0 4
320 400
313 400
313 418
320 418
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
628 692 667 715
640 702 654 717
2 A+
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
635 569 674 592
647 579 661 594
2 B+
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
695 469 734 492
707 479 721 494
2 C+
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
625 342 654 366
635 350 643 366
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
505 344 534 368
515 352 523 368
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
759 87 788 111
769 95 777 111
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
779 95 816 119
789 103 805 119
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
811 106 840 130
821 114 829 130
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
828 127 865 151
838 135 854 151
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
855 148 884 172
865 156 873 172
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
880 166 917 190
890 174 906 190
2 C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
363 347 392 371
373 355 381 371
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
