CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 266 123 0 1 11
0 6
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 M4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4978 0 0
2
43736.5 0
0
13 Logic Switch~
5 220 121 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 M3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9207 0 0
2
43736.5 0
0
13 Logic Switch~
5 168 123 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 M2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6998 0 0
2
43736.5 0
0
13 Logic Switch~
5 116 126 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 M1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3175 0 0
2
43736.5 0
0
14 Logic Display~
6 457 572 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3378 0 0
2
43736.5 0
0
5 4081~
219 414 433 0 3 22
0 5 4 15
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 2 2 0
1 U
922 0 0
2
43736.5 0
0
10 2-In NAND~
219 328 423 0 3 22
0 2 3 5
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6891 0 0
2
43736.5 0
0
10 2-In NAND~
219 318 302 0 3 22
0 11 12 8
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5407 0 0
2
43736.5 0
0
10 2-In NAND~
219 317 251 0 3 22
0 13 11 9
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7349 0 0
2
43736.5 0
0
10 2-In NAND~
219 316 199 0 3 22
0 13 12 10
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3919 0 0
2
43736.5 0
0
5 4023~
219 412 251 0 4 22
0 10 9 8 7
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 3 0
1 U
9747 0 0
2
43736.5 0
0
5 4081~
219 498 334 0 3 22
0 7 6 16
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 1 2 0
1 U
5310 0 0
2
43736.5 0
0
9 Inverter~
13 247 160 0 2 22
0 6 14
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4318 0 0
2
43736.5 0
0
9 Inverter~
13 200 161 0 2 22
0 4 12
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3917 0 0
2
43736.5 0
0
9 Inverter~
13 148 163 0 2 22
0 3 11
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7930 0 0
2
43736.5 0
0
9 Inverter~
13 95 163 0 2 22
0 2 13
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6128 0 0
2
43736.5 0
0
14 Logic Display~
6 457 502 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7346 0 0
2
43736.5 0
0
29
1 0 0 0 0 0 0 9 0 0 3 2
293 242
98 242
1 0 0 0 0 0 0 10 0 0 3 2
292 190
98 190
2 0 0 0 0 0 0 16 0 0 0 2
98 181
98 631
1 0 2 0 0 4096 0 5 0 0 29 2
457 590
116 590
1 0 3 0 0 8192 0 17 0 0 28 3
457 520
457 518
168 518
2 0 4 0 0 4096 0 6 0 0 27 2
390 442
220 442
3 1 5 0 0 8320 0 7 6 0 0 3
355 423
355 424
390 424
2 0 3 0 0 0 0 7 0 0 28 2
304 432
168 432
1 0 2 0 0 0 0 7 0 0 29 2
304 414
116 414
2 0 6 0 0 4096 0 12 0 0 26 2
474 343
266 343
4 1 7 0 0 8320 0 11 12 0 0 4
439 251
454 251
454 325
474 325
3 3 8 0 0 8320 0 8 11 0 0 4
345 302
370 302
370 260
388 260
3 2 9 0 0 4224 0 9 11 0 0 2
344 251
388 251
3 1 10 0 0 8320 0 10 11 0 0 4
343 199
370 199
370 242
388 242
2 0 11 0 0 4096 0 9 0 0 19 2
293 260
151 260
2 0 12 0 0 4096 0 8 0 0 20 2
294 311
203 311
1 0 11 0 0 4096 0 8 0 0 19 2
294 293
151 293
2 0 12 0 0 0 0 10 0 0 20 2
292 208
203 208
2 0 11 0 0 4224 0 15 0 0 0 2
151 181
151 632
2 0 12 0 0 4224 0 14 0 0 0 2
203 179
203 632
2 0 14 0 0 4224 0 13 0 0 0 2
250 178
250 631
1 0 6 0 0 0 0 13 0 0 26 2
250 142
266 142
1 0 4 0 0 0 0 14 0 0 27 2
203 143
220 143
1 0 3 0 0 0 0 15 0 0 28 2
151 145
168 145
1 0 2 0 0 0 0 16 0 0 29 2
98 145
116 145
1 0 6 0 0 4224 0 1 0 0 0 2
266 135
266 630
1 0 4 0 0 4224 0 2 0 0 0 2
220 133
220 630
1 0 3 0 0 4224 0 3 0 0 0 2
168 135
168 631
1 0 2 0 0 4224 0 4 0 0 0 2
116 138
116 632
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
412 559 449 583
422 567 438 583
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
413 484 450 508
423 492 439 508
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
429 404 466 428
439 412 455 428
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
520 306 557 330
530 314 546 330
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
114 48 239 72
124 56 228 72
13 Quest�o 2 TS1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
