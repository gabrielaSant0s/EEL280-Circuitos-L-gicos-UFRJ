CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
90
13 Logic Switch~
5 126 1596 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-4 21 10 29
1 B
-3 13 4 21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9568 0 0
2
43738.8 0
0
13 Logic Switch~
5 108 1596 0 1 11
0 4
0
0 0 21360 90
2 0V
-5 21 9 29
1 A
-3 13 4 21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7178 0 0
2
43738.8 0
0
13 Logic Switch~
5 227 1572 0 1 11
0 8
0
0 0 21360 90
2 0V
-6 23 8 31
1 D
-2 13 5 21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7982 0 0
2
43738.8 0
0
13 Logic Switch~
5 205 1573 0 1 11
0 9
0
0 0 21360 90
2 0V
-5 21 9 29
1 C
-3 13 4 21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
513 0 0
2
43738.8 0
0
13 Logic Switch~
5 575 1573 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8190 0 0
2
43738.8 2
0
13 Logic Switch~
5 571 1525 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5209 0 0
2
43738.8 1
0
13 Logic Switch~
5 573 1474 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7239 0 0
2
43738.8 0
0
13 Logic Switch~
5 581 1035 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9474 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 627 1033 0 1 11
0 36
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3783 0 0
2
5.8991e-315 5.26354e-315
0
13 Logic Switch~
5 665 1033 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 C5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5422 0 0
2
5.8991e-315 5.30499e-315
0
13 Logic Switch~
5 708 1032 0 1 11
0 39
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 D3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8527 0 0
2
5.8991e-315 5.32571e-315
0
13 Logic Switch~
5 234 1016 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
761 0 0
2
5.8991e-315 5.34643e-315
0
13 Logic Switch~
5 191 1017 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 C2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7323 0 0
2
5.8991e-315 5.3568e-315
0
13 Logic Switch~
5 153 1017 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8543 0 0
2
5.8991e-315 5.36716e-315
0
13 Logic Switch~
5 107 1019 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4240 0 0
2
5.8991e-315 5.37752e-315
0
13 Logic Switch~
5 708 463 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7857 0 0
2
43738.8 0
0
13 Logic Switch~
5 665 464 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 C4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7255 0 0
2
43738.8 1
0
13 Logic Switch~
5 627 464 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7736 0 0
2
43738.8 2
0
13 Logic Switch~
5 581 466 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5435 0 0
2
43738.8 3
0
13 Logic Switch~
5 252 477 0 1 11
0 67
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3446 0 0
2
43738.8 4
0
13 Logic Switch~
5 209 478 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 C3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3914 0 0
2
43738.8 5
0
13 Logic Switch~
5 171 478 0 1 11
0 63
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3948 0 0
2
43738.8 6
0
13 Logic Switch~
5 125 480 0 1 11
0 68
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3901 0 0
2
43738.8 7
0
13 Logic Switch~
5 516 110 0 10 11
0 71 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6295 0 0
2
43738.8 8
0
13 Logic Switch~
5 562 109 0 10 11
0 70 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
332 0 0
2
43738.8 9
0
13 Logic Switch~
5 600 109 0 10 11
0 69 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 C1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9737 0 0
2
43738.8 10
0
13 Logic Switch~
5 213 117 0 1 11
0 81
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9910 0 0
2
43738.8 11
0
13 Logic Switch~
5 175 117 0 10 11
0 82 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3834 0 0
2
43738.8 12
0
13 Logic Switch~
5 129 118 0 10 11
0 83 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3138 0 0
2
43738.8 13
0
14 Logic Display~
6 372 1449 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5409 0 0
2
43738.8 0
0
9 Inverter~
13 173 1476 0 2 22
0 7 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U11E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 11 0
1 U
983 0 0
2
43738.8 0
0
9 2-In XOR~
219 115 1541 0 3 22
0 4 3 7
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U23A
27 -3 55 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
6652 0 0
2
43738.8 0
0
7 Ground~
168 371 1396 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4281 0 0
2
43738.8 0
0
7 74LS153
119 277 1485 0 14 29
0 7 6 7 6 9 8 84 85 86
87 2 88 5 89
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
3 U22
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 0 0 0 0
1 U
6847 0 0
2
43738.8 0
0
14 Logic Display~
6 892 1474 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6543 0 0
2
43738.8 0
0
6 74266~
219 819 1505 0 3 22
0 12 11 10
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7168 0 0
2
43738.8 6
0
9 2-In XOR~
219 696 1496 0 3 22
0 14 13 12
0
0 0 624 0
7 74LS386
-24 -24 25 -16
4 U21A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
3828 0 0
2
43738.8 5
0
14 Logic Display~
6 902 642 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
955 0 0
2
43738.8 14
0
5 7413~
219 766 805 0 5 22
0 18 17 16 16 26
0
0 0 624 0
6 74LS13
-14 -24 28 -16
4 U20B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 19 0
1 U
7782 0 0
2
43738.8 15
0
5 7413~
219 766 758 0 5 22
0 17 16 19 19 24
0
0 0 624 0
6 74LS13
-14 -24 28 -16
4 U20A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 19 0
1 U
824 0 0
2
43738.8 16
0
5 7413~
219 766 711 0 5 22
0 22 21 20 20 25
0
0 0 624 0
6 74LS13
-14 -24 28 -16
4 U19B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 18 0
1 U
6983 0 0
2
43738.8 17
0
5 7413~
219 765 659 0 5 22
0 22 23 20 20 27
0
0 0 624 0
6 74LS13
-14 -24 28 -16
4 U19A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 18 0
1 U
3185 0 0
2
43738.8 18
0
5 4011~
219 762 606 0 3 22
0 18 19 28
0
0 0 624 0
4 4011
-7 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 17 0
1 U
4213 0 0
2
43738.8 19
0
5 4011~
219 762 552 0 3 22
0 23 21 29
0
0 0 624 0
4 4011
-7 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 17 0
1 U
9765 0 0
2
43738.8 20
0
10 8-In NAND~
219 865 664 0 9 19
0 29 28 27 25 24 26 24 25 15
0
0 0 624 0
5 74F30
-18 -24 17 -16
3 U17
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
8986 0 0
2
43738.8 21
0
9 Inverter~
13 552 1074 0 2 22
0 37 33
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
3273 0 0
2
5.8991e-315 5.38788e-315
0
9 Inverter~
13 605 1068 0 2 22
0 36 34
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
5636 0 0
2
5.8991e-315 5.39306e-315
0
9 Inverter~
13 646 1070 0 2 22
0 35 41
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
327 0 0
2
5.8991e-315 5.39824e-315
0
9 Inverter~
13 689 1069 0 2 22
0 39 40
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
9233 0 0
2
5.8991e-315 5.40342e-315
0
5 7422~
219 839 1193 0 5 22
0 37 39 37 38 32
0
0 0 624 0
6 74LS22
-21 -28 21 -20
4 U16A
-15 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 16 0
1 U
3875 0 0
2
5.8991e-315 5.4086e-315
0
6 74266~
219 754 1256 0 3 22
0 36 35 38
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9991 0 0
2
5.8991e-315 5.41378e-315
0
5 7422~
219 764 1124 0 5 22
0 34 33 34 33 31
0
0 0 624 0
6 74LS22
-21 -28 21 -20
4 U16B
-15 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 16 0
1 U
3221 0 0
2
5.8991e-315 5.41896e-315
0
5 7422~
219 900 1136 0 5 22
0 31 32 31 32 30
0
0 0 624 0
6 74LS22
-21 -28 21 -20
4 U15A
-15 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 15 0
1 U
8874 0 0
2
5.8991e-315 5.42414e-315
0
14 Logic Display~
6 952 1112 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7400 0 0
2
5.8991e-315 5.42933e-315
0
9 Inverter~
13 215 1053 0 2 22
0 46 52
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
3623 0 0
2
5.8991e-315 5.43192e-315
0
9 Inverter~
13 172 1054 0 2 22
0 49 50
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
3311 0 0
2
5.8991e-315 5.43451e-315
0
9 Inverter~
13 131 1052 0 2 22
0 48 51
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
5736 0 0
2
5.8991e-315 5.4371e-315
0
9 Inverter~
13 78 1058 0 2 22
0 47 53
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
3143 0 0
2
5.8991e-315 5.43969e-315
0
14 Logic Display~
6 416 1186 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5835 0 0
2
5.8991e-315 5.44228e-315
0
5 4082~
219 294 1136 0 5 22
0 47 51 50 46 45
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
5108 0 0
2
5.8991e-315 5.44487e-315
0
5 4082~
219 295 1222 0 5 22
0 46 49 48 47 44
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U12A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
3320 0 0
2
5.8991e-315 5.44746e-315
0
8 3-In OR~
219 366 1204 0 4 22
0 45 44 43 42
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U13A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 13 0
1 U
523 0 0
2
5.8991e-315 5.45005e-315
0
5 4001~
219 282 1292 0 3 22
0 47 46 43
0
0 0 624 0
4 4001
-14 -24 14 -16
4 U14A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 14 0
1 U
3557 0 0
2
5.8991e-315 5.45264e-315
0
9 Inverter~
13 689 500 0 2 22
0 20 19
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
7246 0 0
2
43738.8 22
0
9 Inverter~
13 646 501 0 2 22
0 16 21
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3916 0 0
2
43738.8 23
0
9 Inverter~
13 605 499 0 2 22
0 17 23
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
614 0 0
2
43738.8 24
0
9 Inverter~
13 552 505 0 2 22
0 18 22
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U9B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
8494 0 0
2
43738.8 25
0
14 Logic Display~
6 497 704 0 1 2
10 54
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
774 0 0
2
43738.8 26
0
5 4082~
219 380 662 0 5 22
0 60 59 58 57 55
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
715 0 0
2
43738.8 27
0
5 4081~
219 443 722 0 3 22
0 55 56 54
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
3281 0 0
2
43738.8 28
0
9 Inverter~
13 233 514 0 2 22
0 67 61
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
3593 0 0
2
43738.8 29
0
9 Inverter~
13 190 515 0 2 22
0 65 62
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
7233 0 0
2
43738.8 30
0
9 Inverter~
13 149 513 0 2 22
0 63 66
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
3410 0 0
2
43738.8 31
0
9 Inverter~
13 96 519 0 2 22
0 68 64
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3616 0 0
2
43738.8 32
0
8 4-In OR~
219 288 814 0 5 22
0 64 63 62 61 56
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
5202 0 0
2
43738.8 33
0
8 4-In OR~
219 290 755 0 5 22
0 64 66 65 61 57
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
9145 0 0
2
43738.8 34
0
8 4-In OR~
219 291 698 0 5 22
0 64 63 65 67 58
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
9815 0 0
2
43738.8 35
0
8 4-In OR~
219 291 640 0 5 22
0 68 66 65 67 59
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
4766 0 0
2
43738.8 36
0
8 4-In OR~
219 292 578 0 5 22
0 68 63 62 67 60
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
8325 0 0
2
43738.8 37
0
14 Logic Display~
6 810 173 0 1 2
10 72
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7196 0 0
2
43738.8 38
0
14 Logic Display~
6 441 232 0 1 2
10 74
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3567 0 0
2
43738.8 39
0
8 2-In OR~
219 396 252 0 3 22
0 78 77 74
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
5877 0 0
2
43738.8 40
0
8 2-In OR~
219 337 315 0 3 22
0 76 75 77
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4785 0 0
2
43738.8 41
0
6 74266~
219 659 243 0 3 22
0 70 69 73
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3822 0 0
2
43738.8 42
0
8 2-In OR~
219 755 195 0 3 22
0 71 73 72
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7640 0 0
2
43738.8 43
0
8 2-In OR~
219 332 207 0 3 22
0 80 79 78
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9221 0 0
2
43738.8 44
0
9 2-In AND~
219 264 291 0 3 22
0 82 81 76
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
6484 0 0
2
43738.8 45
0
9 2-In AND~
219 261 172 0 3 22
0 83 82 80
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3689 0 0
2
43738.8 46
0
9 2-In AND~
219 262 229 0 3 22
0 83 81 79
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3952 0 0
2
43738.8 47
0
6 74266~
219 259 357 0 3 22
0 82 81 75
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3631 0 0
2
43738.8 48
0
176
2 1 3 0 0 4224 0 32 1 0 0 2
127 1560
127 1583
1 1 4 0 0 4224 0 32 2 0 0 2
109 1560
109 1583
13 1 5 0 0 4224 0 34 30 0 0 2
309 1467
372 1467
0 2 6 0 0 4096 0 0 34 5 0 3
235 1476
235 1458
245 1458
2 4 6 0 0 4224 0 31 34 0 0 2
194 1476
245 1476
1 0 7 0 0 4096 0 31 0 0 8 2
158 1476
118 1476
0 3 7 0 0 0 0 0 34 8 0 3
232 1449
232 1467
245 1467
3 1 7 0 0 8320 0 32 34 0 0 3
118 1511
118 1449
245 1449
1 6 8 0 0 4224 0 3 34 0 0 3
228 1559
228 1494
245 1494
1 5 9 0 0 4224 0 4 34 0 0 3
206 1560
206 1485
245 1485
1 11 2 0 0 8320 0 33 34 0 0 4
371 1390
325 1390
325 1449
315 1449
3 1 10 0 0 4224 0 36 35 0 0 3
858 1505
892 1505
892 1492
1 2 11 0 0 4224 0 5 36 0 0 4
587 1573
749 1573
749 1514
803 1514
3 1 12 0 0 4224 0 37 36 0 0 2
729 1496
803 1496
1 2 13 0 0 4224 0 6 37 0 0 4
583 1525
638 1525
638 1505
680 1505
1 1 14 0 0 4224 0 7 37 0 0 4
585 1474
643 1474
643 1487
680 1487
9 1 15 0 0 4224 0 45 38 0 0 3
892 664
902 664
902 660
0 9 15 0 0 0 0 0 45 0 0 3
889 667
892 667
892 664
4 0 16 0 0 4096 0 39 0 0 20 3
742 819
733 819
733 810
3 0 16 0 0 4096 0 39 0 0 109 2
742 810
665 810
2 0 17 0 0 4096 0 39 0 0 110 2
742 801
627 801
1 0 18 0 0 4096 0 39 0 0 111 2
742 792
581 792
4 0 19 0 0 4096 0 40 0 0 24 3
742 772
731 772
731 763
3 0 19 0 0 4096 0 40 0 0 100 2
742 763
692 763
2 0 16 0 0 0 0 40 0 0 109 2
742 754
665 754
1 0 17 0 0 0 0 40 0 0 110 2
742 745
627 745
4 0 20 0 0 4096 0 41 0 0 28 3
742 725
732 725
732 716
3 0 20 0 0 4096 0 41 0 0 102 2
742 716
708 716
2 0 21 0 0 4096 0 41 0 0 103 2
742 707
649 707
1 0 22 0 0 4096 0 41 0 0 105 2
742 698
555 698
4 0 20 0 0 0 0 42 0 0 32 3
741 673
732 673
732 664
3 0 20 0 0 0 0 42 0 0 102 2
741 664
708 664
2 0 23 0 0 4096 0 42 0 0 104 2
741 655
608 655
1 0 22 0 0 0 0 42 0 0 105 2
741 646
555 646
2 0 19 0 0 0 0 43 0 0 100 2
738 615
692 615
1 0 18 0 0 0 0 43 0 0 111 2
738 597
581 597
2 0 21 0 0 0 0 44 0 0 103 2
738 561
649 561
1 0 23 0 0 0 0 44 0 0 104 2
738 543
608 543
7 0 24 0 0 4096 0 45 0 0 42 2
841 687
828 687
8 0 25 0 0 8192 0 45 0 0 43 3
841 696
841 698
833 698
5 6 26 0 0 8320 0 39 45 0 0 4
793 805
823 805
823 678
841 678
5 5 24 0 0 8320 0 40 45 0 0 4
793 758
828 758
828 669
841 669
5 4 25 0 0 8320 0 41 45 0 0 4
793 711
833 711
833 660
841 660
5 3 27 0 0 4224 0 42 45 0 0 4
792 659
833 659
833 651
841 651
3 2 28 0 0 4224 0 43 45 0 0 4
789 606
828 606
828 642
841 642
3 1 29 0 0 8320 0 44 45 0 0 4
789 552
833 552
833 633
841 633
5 1 30 0 0 4224 0 53 54 0 0 3
927 1136
952 1136
952 1130
1 0 31 0 0 4096 0 53 0 0 51 3
876 1118
865 1118
865 1124
4 0 32 0 0 4096 0 53 0 0 50 2
876 1154
870 1154
5 2 32 0 0 8320 0 50 53 0 0 4
866 1193
870 1193
870 1142
876 1142
5 3 31 0 0 4224 0 52 53 0 0 4
791 1124
868 1124
868 1130
876 1130
4 0 33 0 0 8192 0 52 0 0 55 3
740 1142
732 1142
732 1130
1 0 34 0 0 8192 0 52 0 0 54 3
740 1106
732 1106
732 1118
3 0 34 0 0 4096 0 52 0 0 70 2
740 1118
608 1118
2 0 33 0 0 4096 0 52 0 0 71 2
740 1130
555 1130
2 0 35 0 0 4096 0 51 0 0 64 2
738 1265
665 1265
1 0 36 0 0 4096 0 51 0 0 65 2
738 1247
627 1247
1 0 37 0 0 4096 0 50 0 0 61 3
815 1175
796 1175
796 1187
3 4 38 0 0 4224 0 51 50 0 0 3
793 1256
793 1211
815 1211
2 0 39 0 0 4096 0 50 0 0 68 2
815 1199
708 1199
3 0 37 0 0 4096 0 50 0 0 73 2
815 1187
581 1187
1 0 35 0 0 0 0 48 0 0 64 2
649 1052
665 1052
1 0 36 0 0 0 0 47 0 0 65 2
608 1050
627 1050
1 0 35 0 0 4224 0 10 0 0 0 2
665 1045
665 1291
1 0 36 0 0 4224 0 9 0 0 0 2
627 1045
627 1292
2 0 40 0 0 4224 0 49 0 0 0 2
692 1087
692 1291
1 0 39 0 0 0 0 49 0 0 68 2
692 1051
708 1051
1 0 39 0 0 4224 0 11 0 0 0 2
708 1044
708 1289
2 0 41 0 0 4224 0 48 0 0 0 2
649 1088
649 1289
2 0 34 0 0 4224 0 47 0 0 0 2
608 1086
608 1293
2 0 33 0 0 4224 0 46 0 0 0 2
555 1092
555 1293
1 0 37 0 0 0 0 46 0 0 73 2
555 1056
581 1056
1 0 37 0 0 4224 0 8 0 0 0 2
581 1047
581 1293
4 1 42 0 0 4224 0 62 59 0 0 2
399 1204
416 1204
3 3 43 0 0 8320 0 63 62 0 0 4
321 1292
340 1292
340 1213
353 1213
5 2 44 0 0 4224 0 61 62 0 0 4
316 1222
345 1222
345 1204
354 1204
5 1 45 0 0 8320 0 60 62 0 0 4
315 1136
345 1136
345 1195
353 1195
2 0 46 0 0 4096 0 63 0 0 94 2
269 1301
234 1301
1 0 47 0 0 4096 0 63 0 0 99 2
269 1283
107 1283
1 0 46 0 0 4096 0 61 0 0 94 2
271 1209
234 1209
4 0 47 0 0 4096 0 61 0 0 99 2
271 1236
107 1236
3 0 48 0 0 4096 0 61 0 0 91 2
271 1227
153 1227
2 0 49 0 0 4096 0 61 0 0 90 2
271 1218
191 1218
4 0 46 0 0 0 0 60 0 0 94 2
270 1150
234 1150
3 0 50 0 0 4096 0 60 0 0 95 2
270 1141
175 1141
2 0 51 0 0 4096 0 60 0 0 96 2
270 1132
134 1132
1 0 47 0 0 0 0 60 0 0 99 2
270 1123
107 1123
1 0 48 0 0 0 0 57 0 0 91 2
134 1034
153 1034
1 0 49 0 0 0 0 56 0 0 90 2
175 1036
191 1036
1 0 49 0 0 4224 0 13 0 0 0 2
191 1029
191 1330
1 0 48 0 0 4224 0 14 0 0 0 2
153 1029
153 1330
2 0 52 0 0 4224 0 55 0 0 0 2
218 1071
218 1329
1 0 46 0 0 0 0 55 0 0 94 2
218 1035
234 1035
1 0 46 0 0 4224 0 12 0 0 0 2
234 1028
234 1328
2 0 50 0 0 4224 0 56 0 0 0 2
175 1072
175 1330
2 0 51 0 0 4224 0 57 0 0 0 2
134 1070
134 1331
2 0 53 0 0 4224 0 58 0 0 0 2
81 1076
81 1330
1 0 47 0 0 0 0 58 0 0 99 2
81 1040
107 1040
1 0 47 0 0 4224 0 15 0 0 0 2
107 1031
107 1332
2 0 19 0 0 4224 0 64 0 0 0 2
692 518
692 863
1 0 20 0 0 0 0 64 0 0 102 2
692 482
708 482
1 0 20 0 0 4224 0 16 0 0 0 2
708 475
708 864
2 0 21 0 0 4224 0 65 0 0 0 2
649 519
649 864
2 0 23 0 0 4224 0 66 0 0 0 2
608 517
608 863
2 0 22 0 0 4224 0 67 0 0 0 2
555 523
555 867
1 0 18 0 0 0 0 67 0 0 111 2
555 487
581 487
1 0 16 0 0 0 0 65 0 0 109 2
649 483
665 483
1 0 17 0 0 0 0 66 0 0 110 2
608 481
627 481
1 0 16 0 0 4224 0 17 0 0 0 2
665 476
665 865
1 0 17 0 0 4224 0 18 0 0 0 2
627 476
627 866
1 0 18 0 0 4224 0 19 0 0 0 2
581 478
581 867
3 1 54 0 0 4224 0 70 68 0 0 2
464 722
497 722
5 1 55 0 0 8320 0 69 70 0 0 4
401 662
405 662
405 713
419 713
5 2 56 0 0 8320 0 75 70 0 0 4
321 814
397 814
397 731
419 731
5 4 57 0 0 8320 0 76 69 0 0 4
323 755
343 755
343 676
356 676
5 3 58 0 0 8320 0 77 69 0 0 4
324 698
348 698
348 667
356 667
5 2 59 0 0 4224 0 78 69 0 0 4
324 640
343 640
343 658
356 658
5 1 60 0 0 8320 0 79 69 0 0 4
325 578
348 578
348 649
356 649
4 0 61 0 0 4096 0 75 0 0 139 2
271 828
236 828
3 0 62 0 0 4096 0 75 0 0 142 2
271 819
193 819
2 0 63 0 0 4096 0 75 0 0 149 2
271 810
171 810
1 0 64 0 0 4096 0 75 0 0 144 2
271 801
99 801
4 0 61 0 0 4096 0 76 0 0 139 2
273 769
236 769
3 0 65 0 0 4096 0 76 0 0 148 2
273 760
209 760
2 0 66 0 0 4096 0 76 0 0 143 2
273 751
152 751
1 0 64 0 0 4096 0 76 0 0 144 2
273 742
99 742
4 0 67 0 0 4096 0 77 0 0 141 2
274 712
252 712
3 0 65 0 0 4096 0 77 0 0 148 2
274 703
209 703
2 0 63 0 0 4096 0 77 0 0 149 2
274 694
171 694
1 0 64 0 0 4096 0 77 0 0 144 2
274 685
99 685
4 0 67 0 0 0 0 78 0 0 141 2
274 654
252 654
3 0 65 0 0 0 0 78 0 0 148 2
274 645
209 645
2 0 66 0 0 4096 0 78 0 0 143 2
274 636
152 636
1 0 68 0 0 4096 0 78 0 0 150 2
274 627
125 627
4 0 67 0 0 4096 0 79 0 0 141 2
275 592
252 592
3 0 62 0 0 4096 0 79 0 0 142 2
275 583
193 583
2 0 63 0 0 4096 0 79 0 0 149 2
275 574
171 574
1 0 68 0 0 4096 0 79 0 0 150 2
275 565
125 565
2 0 61 0 0 4224 0 71 0 0 0 2
236 532
236 877
1 0 67 0 0 0 0 71 0 0 141 2
236 496
252 496
1 0 67 0 0 4224 0 20 0 0 0 2
252 489
252 878
2 0 62 0 0 4224 0 72 0 0 0 2
193 533
193 878
2 0 66 0 0 4224 0 73 0 0 0 2
152 531
152 877
2 0 64 0 0 4224 0 74 0 0 0 2
99 537
99 881
1 0 68 0 0 0 0 74 0 0 150 2
99 501
125 501
1 0 65 0 0 0 0 72 0 0 148 2
193 497
209 497
1 0 63 0 0 0 0 73 0 0 149 2
152 495
171 495
1 0 65 0 0 4224 0 21 0 0 0 2
209 490
209 879
1 0 63 0 0 4224 0 22 0 0 0 2
171 490
171 880
1 0 68 0 0 4224 0 23 0 0 0 2
125 492
125 881
2 0 69 0 0 4096 0 84 0 0 171 2
643 252
600 252
1 0 70 0 0 4096 0 84 0 0 172 2
643 234
562 234
1 0 71 0 0 4224 0 85 0 0 173 2
742 186
516 186
3 1 72 0 0 4224 0 85 80 0 0 3
788 195
810 195
810 191
3 2 73 0 0 8320 0 84 85 0 0 4
698 243
734 243
734 204
742 204
3 1 74 0 0 8320 0 82 81 0 0 3
429 252
429 250
441 250
3 2 75 0 0 8320 0 90 83 0 0 4
298 357
316 357
316 324
324 324
3 1 76 0 0 4224 0 87 83 0 0 4
285 291
316 291
316 306
324 306
3 2 77 0 0 8320 0 83 82 0 0 4
370 315
375 315
375 261
383 261
3 1 78 0 0 8320 0 86 82 0 0 4
365 207
375 207
375 243
383 243
3 2 79 0 0 12416 0 89 86 0 0 4
283 229
289 229
289 216
319 216
3 1 80 0 0 8320 0 88 86 0 0 3
282 172
282 198
319 198
2 0 81 0 0 4096 0 90 0 0 174 2
243 366
213 366
1 0 82 0 0 4096 0 90 0 0 175 2
243 348
175 348
2 0 81 0 0 0 0 87 0 0 174 2
240 300
213 300
1 0 82 0 0 0 0 87 0 0 175 2
240 282
175 282
2 0 81 0 0 0 0 89 0 0 174 2
238 238
213 238
1 0 83 0 0 4096 0 89 0 0 176 2
238 220
129 220
2 0 82 0 0 0 0 88 0 0 175 2
237 181
175 181
1 0 83 0 0 0 0 88 0 0 176 2
237 163
129 163
1 0 69 0 0 4224 0 26 0 0 0 2
600 121
600 315
1 0 70 0 0 4224 0 25 0 0 0 2
562 121
562 316
1 0 71 0 0 0 0 24 0 0 0 2
516 122
516 314
1 0 81 0 0 4224 0 27 0 0 0 2
213 129
213 400
1 0 82 0 0 4224 0 28 0 0 0 2
175 129
175 397
1 0 83 0 0 4224 0 29 0 0 0 2
129 130
129 401
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
70 1378 251 1402
80 1386 240 1402
20 LETRA D N�O REDUZIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
594 1375 743 1399
604 1383 732 1399
16 LETRA D REDUZIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
782 1379 931 1403
792 1387 920 1403
16 D xnor (A xor B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
571 397 720 421
581 405 709 421
16 LETRA B REDUZIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
106 406 287 430
116 414 276 430
20 LETRA B NAO REDUZIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
493 31 714 55
503 39 703 55
25 LETRA A NUMERO 1 REDUZIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
111 33 364 57
121 41 353 57
29 LETRA A NUMERO 1 NAO REDUZIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
87 941 268 965
97 949 257 965
20 LETRA C NAO REDUZIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
569 945 718 969
579 953 707 969
16 LETRA C REDUZIDA
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
