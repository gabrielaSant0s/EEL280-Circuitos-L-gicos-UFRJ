CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 662 261 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3641 0 0
2
43727.1 4
0
13 Logic Switch~
5 662 303 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3104 0 0
2
43727.1 3
0
5 4030~
219 765 270 0 3 22
0 14 13 15
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3296 0 0
2
43727.1 2
0
7 Ground~
168 901 356 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8534 0 0
2
43727.1 1
0
4 LED~
171 901 318 0 1 2
10 15
0
0 0 880 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
949 0 0
2
43727.1 0
0
4 LED~
171 961 136 0 1 2
10 16
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3371 0 0
2
43727.1 8
0
7 Ground~
168 961 160 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7311 0 0
2
43727.1 7
0
5 4011~
219 908 125 0 3 22
0 18 17 16
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 9 0
1 U
3409 0 0
2
43727.1 6
0
5 4011~
219 833 167 0 3 22
0 14 19 18
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 8 0
1 U
3526 0 0
2
43727.1 5
0
5 4011~
219 760 137 0 3 22
0 14 13 19
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 8 0
1 U
4129 0 0
2
43727.1 4
0
5 4011~
219 757 83 0 3 22
0 14 13 19
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 8 0
1 U
6278 0 0
2
43727.1 3
0
5 4011~
219 836 92 0 3 22
0 14 19 18
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 8 0
1 U
3482 0 0
2
43727.1 2
0
13 Logic Switch~
5 657 74 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8323 0 0
2
43727.1 1
0
13 Logic Switch~
5 658 129 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3984 0 0
2
43727.1 0
0
13 Logic Switch~
5 582 670 0 1 11
0 7
0
0 0 21344 0
2 0V
-8 -16 6 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7622 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 583 632 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
816 0 0
2
5.89908e-315 5.26354e-315
0
13 Logic Switch~
5 581 593 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4656 0 0
2
5.89908e-315 5.30499e-315
0
13 Logic Switch~
5 581 551 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6356 0 0
2
5.89908e-315 5.32571e-315
0
13 Logic Switch~
5 583 516 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7479 0 0
2
5.89908e-315 5.34643e-315
0
13 Logic Switch~
5 584 471 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5690 0 0
2
5.89908e-315 5.3568e-315
0
4 LED~
171 924 583 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5617 0 0
2
5.89908e-315 5.36716e-315
0
7 Ground~
168 924 610 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3903 0 0
2
5.89908e-315 5.37752e-315
0
5 4073~
219 844 560 0 4 22
0 4 5 6 3
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
4452 0 0
2
5.89908e-315 5.38788e-315
0
10 2-In XNOR~
219 722 647 0 3 22
0 8 7 6
0
0 0 608 0
4 4077
-7 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
6282 0 0
2
5.89908e-315 5.39306e-315
0
10 2-In XNOR~
219 722 569 0 3 22
0 10 9 5
0
0 0 608 0
4 4077
-7 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
7187 0 0
2
5.89908e-315 5.39824e-315
0
10 2-In XNOR~
219 719 493 0 3 22
0 12 11 4
0
0 0 608 0
4 4077
-7 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
6866 0 0
2
5.89908e-315 5.40342e-315
0
27
1 2 0 0 0 0 0 2 3 0 0 4
674 303
700 303
700 279
749 279
1 1 0 0 0 0 0 3 1 0 0 2
749 261
674 261
2 1 2 0 0 0 0 5 4 0 0 2
901 328
901 350
3 1 15 0 0 0 0 3 5 0 0 3
798 270
901 270
901 308
3 2 0 0 0 0 0 10 12 0 0 4
787 137
799 137
799 101
812 101
3 1 0 0 0 0 0 12 8 0 0 3
863 92
863 116
884 116
3 2 0 0 0 0 0 9 8 0 0 4
860 167
873 167
873 134
884 134
2 1 2 0 0 0 0 6 7 0 0 2
961 146
961 154
3 1 16 0 0 0 0 8 6 0 0 4
935 125
949 125
949 126
961 126
0 2 0 0 0 0 0 0 9 14 0 3
676 129
676 176
809 176
0 1 0 0 0 0 0 0 9 16 0 5
677 74
677 38
621 38
621 158
809 158
3 1 0 0 0 0 0 11 12 0 0 2
784 83
812 83
2 0 0 0 0 0 0 10 0 0 14 3
736 146
690 146
690 129
1 1 0 0 0 0 0 10 14 0 0 4
736 128
690 128
690 129
670 129
2 0 0 0 0 0 0 11 0 0 16 3
733 92
689 92
689 74
1 1 0 0 0 0 0 13 11 0 0 2
669 74
733 74
1 2 2 0 0 4096 0 22 21 0 0 2
924 604
924 593
4 1 3 0 0 4224 0 23 21 0 0 3
865 560
924 560
924 573
3 1 4 0 0 8320 0 26 23 0 0 4
758 493
812 493
812 551
820 551
3 2 5 0 0 4224 0 25 23 0 0 4
761 569
807 569
807 560
820 560
3 3 6 0 0 8320 0 24 23 0 0 4
761 647
812 647
812 569
820 569
1 2 7 0 0 12416 0 15 24 0 0 4
594 670
637 670
637 656
706 656
1 1 8 0 0 8320 0 18 24 0 0 4
593 551
637 551
637 638
706 638
1 2 9 0 0 4224 0 16 25 0 0 4
595 632
671 632
671 578
706 578
1 1 10 0 0 4224 0 19 25 0 0 4
595 516
671 516
671 560
706 560
1 2 11 0 0 4224 0 17 26 0 0 4
593 593
696 593
696 502
703 502
1 1 12 0 0 4224 0 20 26 0 0 4
596 471
695 471
695 484
703 484
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 127
80 367 1117 391
90 375 1106 391
127 #------------------------------------------------------------------------------------------------------------------------------
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 78
133 427 266 551
143 435 255 531
78 A B | A XNor B 
 
0 0 |   1     
0 1 |   0     
1 0 |   0     
1 1 |   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
136 382 245 406
146 390 234 406
11 Quest�o 4 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
694 213 875 237
704 221 864 237
20 F = A'B'+AB com XNOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
653 7 906 31
663 15 895 31
29 F = A'B' + AB com portas NAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
130 70 255 94
140 78 244 94
13 F = A'B' + AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 124
132 114 409 218
142 122 398 202
124 A B | A . B | A'. B'| A'.B'+ A.B
0 0 |   0   |	1   |	1
0 1 |   0   |	0   |	0
1 0 |   0   |	0   |	0
1 1 |   1   |	0   |	1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
126 24 235 48
136 32 224 48
11 Quest�o 4 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 154
125 547 482 691
135 555 471 667
154 bits  : A = A2,A1,A0
	B = B2,B1,B0

C = (A2 Nxor B2).(A1 Nxor B1).(A0 Nxor B0)

Se C = 1 ent�o A e B s�o iguais 
Se C = 0 ent�o A e B s�o diferentes
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
