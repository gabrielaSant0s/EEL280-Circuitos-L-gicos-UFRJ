CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
530 460 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.168350
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
58
13 Logic Switch~
5 729 1474 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Rbi
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 1105 530 0 1 11
0 29
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 LT
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 429 279 0 1 11
0 35
0
0 0 21360 270
2 0V
-7 -21 7 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89909e-315 5.32571e-315
0
13 Logic Switch~
5 486 276 0 1 11
0 32
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89909e-315 5.30499e-315
0
13 Logic Switch~
5 538 276 0 1 11
0 30
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 W
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89909e-315 5.26354e-315
0
13 Logic Switch~
5 602 278 0 1 11
0 47
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89909e-315 0
0
2 +V
167 733 1601 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8901 0 0
2
5.89909e-315 0
0
5 4082~
219 660 1513 0 5 22
0 34 33 31 57 4
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U23A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 25 0
1 U
7361 0 0
2
5.89909e-315 0
0
9 Inverter~
13 774 1474 0 2 22
0 5 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
4747 0 0
2
5.89909e-315 0
0
10 3-In NAND~
219 840 1513 0 4 22
0 6 4 3 7
0
0 0 624 0
6 74LS10
-21 -28 21 -20
4 U22A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 24 0
1 U
972 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 1019 1311 0 3 22
0 21 7 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U21D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 23 0
1 U
3472 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 1015 1129 0 3 22
0 19 7 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U21C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 23 0
1 U
9998 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 1017 986 0 3 22
0 17 7 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U21B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 23 0
1 U
3536 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 1017 794 0 3 22
0 16 7 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 23 0
1 U
4597 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 1018 624 0 3 22
0 15 7 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 20 0
1 U
3835 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 1018 541 0 3 22
0 14 7 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
3670 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 1018 459 0 3 22
0 9 7 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
5616 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 1159 1309 0 3 22
0 20 29 22
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 22 0
1 U
9323 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 1160 1182 0 3 22
0 18 29 23
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
317 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 1155 1065 0 3 22
0 13 29 24
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U16A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
3108 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 1149 957 0 3 22
0 11 29 25
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 1146 863 0 3 22
0 12 29 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 21 0
1 U
9672 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 1144 766 0 3 22
0 10 29 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 21 0
1 U
7876 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 1143 670 0 3 22
0 8 29 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
6369 0 0
2
5.89909e-315 0
0
14 Logic Display~
6 1105 1435 0 1 2
10 29
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89909e-315 0
0
9 Inverter~
13 394 361 0 2 22
0 35 57
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
7100 0 0
2
5.89909e-315 5.47595e-315
0
9 Inverter~
13 455 360 0 2 22
0 32 31
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3820 0 0
2
5.89909e-315 5.47466e-315
0
9 Inverter~
13 511 363 0 2 22
0 30 33
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
7678 0 0
2
5.89909e-315 5.47336e-315
0
9 Inverter~
13 572 365 0 2 22
0 47 34
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
961 0 0
2
5.89909e-315 5.47207e-315
0
6 74266~
219 702 493 0 3 22
0 32 47 55
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3178 0 0
2
5.89909e-315 5.47077e-315
0
8 2-In OR~
219 797 450 0 3 22
0 56 55 9
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3409 0 0
2
5.89909e-315 5.46818e-315
0
8 2-In OR~
219 700 417 0 3 22
0 35 30 56
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3951 0 0
2
5.89909e-315 5.46559e-315
0
8 2-In OR~
219 803 532 0 3 22
0 31 54 14
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8885 0 0
2
5.89909e-315 5.463e-315
0
6 74266~
219 681 581 0 3 22
0 30 47 54
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3780 0 0
2
5.89909e-315 5.46041e-315
0
8 2-In OR~
219 724 640 0 3 22
0 33 47 53
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
9265 0 0
2
5.89909e-315 5.45782e-315
0
8 2-In OR~
219 807 614 0 3 22
0 32 53 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
9442 0 0
2
5.89909e-315 5.45523e-315
0
9 2-In AND~
219 709 817 0 3 22
0 31 30 51
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
9424 0 0
2
5.89909e-315 5.45264e-315
0
9 2-In AND~
219 714 759 0 3 22
0 31 34 48
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
9968 0 0
2
5.89909e-315 5.45005e-315
0
9 2-In AND~
219 715 710 0 3 22
0 34 30 49
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
9281 0 0
2
5.89909e-315 5.44746e-315
0
8 3-In OR~
219 797 699 0 4 22
0 35 49 48 52
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
8464 0 0
2
5.89909e-315 5.44487e-315
0
8 3-In OR~
219 868 782 0 4 22
0 52 51 50 16
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
7168 0 0
2
5.89909e-315 5.44228e-315
0
9 3-In AND~
219 711 865 0 4 22
0 33 47 32 50
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 6 0
1 U
3171 0 0
2
5.89909e-315 5.43969e-315
0
8 2-In OR~
219 758 946 0 3 22
0 31 30 46
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
4139 0 0
2
5.89909e-315 5.4371e-315
0
9 2-In AND~
219 865 975 0 3 22
0 46 34 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6435 0 0
2
5.89909e-315 5.43451e-315
0
9 2-In AND~
219 717 1187 0 3 22
0 33 34 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
5283 0 0
2
5.89909e-315 5.43192e-315
0
9 2-In AND~
219 720 1128 0 3 22
0 32 33 44
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
6874 0 0
2
5.89909e-315 5.42933e-315
0
9 2-In AND~
219 721 1061 0 3 22
0 32 34 45
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
5305 0 0
2
5.89909e-315 5.42414e-315
0
8 2-In OR~
219 797 1084 0 3 22
0 45 35 42
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
34 0 0
2
5.89909e-315 5.41896e-315
0
8 2-In OR~
219 794 1159 0 3 22
0 44 43 41
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
969 0 0
2
5.89909e-315 5.41378e-315
0
8 2-In OR~
219 869 1121 0 3 22
0 42 41 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
8402 0 0
2
5.89909e-315 5.4086e-315
0
9 2-In AND~
219 727 1380 0 3 22
0 30 34 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
3751 0 0
2
5.89909e-315 5.40342e-315
0
9 2-In AND~
219 728 1321 0 3 22
0 32 33 39
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
4292 0 0
2
5.89909e-315 5.39824e-315
0
9 2-In AND~
219 728 1263 0 3 22
0 30 31 37
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
6118 0 0
2
5.89909e-315 5.39306e-315
0
8 2-In OR~
219 891 1302 0 3 22
0 40 36 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
34 0 0
2
5.89909e-315 5.38788e-315
0
8 2-In OR~
219 820 1353 0 3 22
0 39 38 36
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
6357 0 0
2
5.89909e-315 5.37752e-315
0
8 2-In OR~
219 827 1242 0 3 22
0 35 37 40
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
319 0 0
2
5.89909e-315 5.36716e-315
0
9 CC 7-Seg~
183 1257 586 0 17 19
10 28 27 26 25 24 23 22 58 2
0 0 0 0 0 0 0 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3976 0 0
2
5.89909e-315 5.3568e-315
0
7 Ground~
168 1357 654 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7634 0 0
2
5.89909e-315 5.34643e-315
0
112
3 1 3 0 0 4224 0 10 7 0 0 3
816 1522
816 1610
733 1610
5 2 4 0 0 4224 0 8 10 0 0 2
681 1513
816 1513
1 1 5 0 0 4224 0 1 9 0 0 2
741 1474
759 1474
1 2 6 0 0 4224 0 10 9 0 0 3
816 1504
816 1474
795 1474
2 0 7 0 0 4096 0 11 0 0 12 2
995 1320
984 1320
2 0 7 0 0 0 0 12 0 0 12 2
991 1138
984 1138
2 0 7 0 0 0 0 13 0 0 12 2
993 995
984 995
2 0 7 0 0 0 0 14 0 0 12 2
993 803
984 803
2 0 7 0 0 0 0 15 0 0 12 2
994 633
984 633
2 0 7 0 0 0 0 16 0 0 12 2
994 550
984 550
2 0 7 0 0 0 0 17 0 0 12 2
994 468
984 468
4 0 7 0 0 8320 0 10 0 0 0 4
867 1513
984 1513
984 334
1007 334
3 1 8 0 0 8320 0 17 24 0 0 4
1039 459
1071 459
1071 661
1130 661
1 3 9 0 0 4224 0 17 31 0 0 2
994 450
830 450
3 1 10 0 0 8320 0 16 23 0 0 4
1039 541
1057 541
1057 757
1131 757
3 1 11 0 0 4224 0 14 21 0 0 3
1038 794
1038 948
1136 948
3 1 12 0 0 8320 0 15 22 0 0 4
1039 624
1044 624
1044 854
1133 854
3 1 13 0 0 8320 0 13 20 0 0 4
1038 986
1078 986
1078 1056
1142 1056
3 1 14 0 0 4224 0 33 16 0 0 2
836 532
994 532
3 1 15 0 0 8320 0 36 15 0 0 3
840 614
840 615
994 615
4 1 16 0 0 8320 0 41 14 0 0 3
901 782
901 785
993 785
3 1 17 0 0 8320 0 44 13 0 0 3
886 975
886 977
993 977
3 1 18 0 0 4224 0 12 19 0 0 4
1036 1129
1121 1129
1121 1173
1147 1173
3 1 19 0 0 8320 0 50 12 0 0 3
902 1121
902 1120
991 1120
3 1 20 0 0 4224 0 11 18 0 0 6
1040 1311
1122 1311
1122 1299
1121 1299
1121 1300
1146 1300
3 1 21 0 0 4224 0 54 11 0 0 2
924 1302
995 1302
7 3 22 0 0 4224 0 57 18 0 0 3
1272 622
1272 1309
1192 1309
6 3 23 0 0 4224 0 57 19 0 0 3
1266 622
1266 1182
1193 1182
5 3 24 0 0 4224 0 57 20 0 0 3
1260 622
1260 1065
1188 1065
4 3 25 0 0 4224 0 57 21 0 0 3
1254 622
1254 957
1182 957
3 3 26 0 0 4224 0 57 22 0 0 3
1248 622
1248 863
1179 863
2 3 27 0 0 4224 0 57 23 0 0 3
1242 622
1242 766
1177 766
1 3 28 0 0 8320 0 57 24 0 0 3
1236 622
1236 670
1176 670
2 0 29 0 0 4096 0 18 0 0 41 2
1146 1318
1105 1318
2 0 29 0 0 4096 0 19 0 0 41 2
1147 1191
1105 1191
2 0 29 0 0 0 0 20 0 0 41 2
1142 1074
1105 1074
2 0 29 0 0 0 0 21 0 0 41 2
1136 966
1105 966
2 0 29 0 0 0 0 22 0 0 41 2
1133 872
1105 872
2 0 29 0 0 0 0 23 0 0 41 2
1131 775
1105 775
2 0 29 0 0 0 0 24 0 0 41 2
1130 679
1105 679
1 1 29 0 0 4224 0 2 25 0 0 2
1105 542
1105 1421
1 9 2 0 0 4224 0 58 57 0 0 4
1357 648
1357 519
1257 519
1257 544
1 0 30 0 0 4096 0 53 0 0 105 2
704 1254
538 1254
2 0 31 0 0 4096 0 53 0 0 108 2
704 1272
458 1272
1 0 32 0 0 4096 0 52 0 0 109 2
704 1312
486 1312
2 0 33 0 0 4096 0 52 0 0 104 2
704 1330
514 1330
2 0 34 0 0 4096 0 51 0 0 102 2
703 1389
575 1389
1 0 30 0 0 0 0 51 0 0 105 2
703 1371
538 1371
1 0 35 0 0 4096 0 56 0 0 112 2
814 1233
428 1233
3 2 36 0 0 8320 0 55 54 0 0 4
853 1353
870 1353
870 1311
878 1311
3 2 37 0 0 4224 0 53 56 0 0 4
749 1263
783 1263
783 1251
814 1251
3 2 38 0 0 4224 0 51 55 0 0 4
748 1380
788 1380
788 1362
807 1362
3 1 39 0 0 4224 0 52 55 0 0 4
749 1321
788 1321
788 1344
807 1344
3 1 40 0 0 4224 0 56 54 0 0 3
860 1242
860 1293
878 1293
2 0 34 0 0 0 0 45 0 0 102 2
693 1196
575 1196
2 0 33 0 0 0 0 46 0 0 104 2
696 1137
514 1137
1 0 33 0 0 0 0 45 0 0 104 2
693 1178
514 1178
2 0 34 0 0 0 0 47 0 0 102 2
697 1070
575 1070
1 0 32 0 0 0 0 47 0 0 109 2
697 1052
486 1052
2 0 35 0 0 0 0 48 0 0 112 2
784 1093
428 1093
3 2 41 0 0 8320 0 49 50 0 0 4
827 1159
848 1159
848 1130
856 1130
3 1 42 0 0 8320 0 48 50 0 0 4
830 1084
848 1084
848 1112
856 1112
3 2 43 0 0 4224 0 45 49 0 0 4
738 1187
773 1187
773 1168
781 1168
3 1 44 0 0 4224 0 46 49 0 0 4
741 1128
773 1128
773 1150
781 1150
3 1 45 0 0 8320 0 47 48 0 0 3
742 1061
742 1075
784 1075
0 1 32 0 0 0 0 0 46 109 0 2
486 1119
696 1119
0 2 34 0 0 4096 0 0 44 102 0 4
575 1010
825 1010
825 984
841 984
3 1 46 0 0 4224 0 43 44 0 0 4
791 946
824 946
824 966
841 966
0 2 30 0 0 4096 0 0 43 105 0 4
538 970
708 970
708 955
745 955
0 1 31 0 0 4096 0 0 43 108 0 4
458 922
708 922
708 937
745 937
3 0 32 0 0 0 0 42 0 0 109 2
687 874
486 874
2 0 47 0 0 4096 0 42 0 0 101 2
687 865
602 865
1 0 33 0 0 0 0 42 0 0 104 2
687 856
514 856
2 0 30 0 0 0 0 37 0 0 105 2
685 826
538 826
1 0 31 0 0 0 0 37 0 0 108 2
685 808
458 808
2 0 34 0 0 0 0 38 0 0 102 2
690 768
575 768
1 0 34 0 0 0 0 39 0 0 102 2
691 701
575 701
1 0 31 0 0 0 0 38 0 0 108 2
690 750
458 750
2 0 30 0 0 0 0 39 0 0 105 2
691 719
538 719
3 3 48 0 0 8320 0 38 40 0 0 4
735 759
764 759
764 708
784 708
3 2 49 0 0 12416 0 39 40 0 0 4
736 710
752 710
752 699
785 699
1 0 35 0 0 0 0 40 0 0 112 2
784 690
428 690
4 3 50 0 0 4224 0 42 41 0 0 4
732 865
832 865
832 791
855 791
3 2 51 0 0 4224 0 37 41 0 0 4
730 817
807 817
807 782
856 782
4 1 52 0 0 8320 0 40 41 0 0 4
830 699
847 699
847 773
855 773
1 0 33 0 0 4096 0 35 0 0 104 2
711 631
514 631
2 0 47 0 0 4096 0 35 0 0 101 2
711 649
602 649
1 0 32 0 0 4096 0 36 0 0 109 2
794 605
486 605
3 2 53 0 0 4224 0 35 36 0 0 4
757 640
786 640
786 623
794 623
2 0 47 0 0 0 0 34 0 0 101 2
665 590
602 590
1 0 30 0 0 0 0 34 0 0 105 2
665 572
538 572
1 0 31 0 0 4096 0 33 0 0 108 2
790 523
458 523
3 2 54 0 0 8320 0 34 33 0 0 3
720 581
720 541
790 541
2 0 47 0 0 0 0 30 0 0 101 2
686 502
602 502
1 0 35 0 0 0 0 32 0 0 112 2
687 408
428 408
3 2 55 0 0 4224 0 30 31 0 0 4
741 493
776 493
776 459
784 459
0 1 32 0 0 0 0 0 30 109 0 4
486 449
679 449
679 484
686 484
0 2 30 0 0 0 0 0 32 105 0 4
538 489
661 489
661 426
687 426
3 1 56 0 0 4224 0 32 31 0 0 4
733 417
764 417
764 441
784 441
0 1 47 0 0 0 0 0 29 101 0 3
602 338
575 338
575 347
1 0 47 0 0 4224 0 6 0 0 0 2
602 290
602 1438
2 1 34 0 0 4224 0 29 8 0 0 3
575 383
575 1500
636 1500
1 0 30 0 0 0 0 28 0 0 105 2
514 345
538 345
2 2 33 0 0 4224 0 28 8 0 0 3
514 381
514 1509
636 1509
1 0 30 0 0 4224 0 5 0 0 0 2
538 288
538 1441
1 0 32 0 0 0 0 27 0 0 109 2
458 342
486 342
1 0 35 0 0 0 0 26 0 0 112 2
397 343
428 343
2 3 31 0 0 4224 0 27 8 0 0 3
458 378
458 1518
636 1518
1 0 32 0 0 4224 0 4 0 0 0 2
486 288
486 1443
1 0 32 0 0 0 0 4 0 0 0 2
486 288
486 885
2 4 57 0 0 4224 0 26 8 0 0 3
397 379
397 1527
636 1527
1 0 35 0 0 12416 0 3 0 0 0 4
429 291
429 343
428 343
428 1445
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
388 188 641 212
398 196 630 212
29 Decodificador BCD 7 segmentos
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
897 728 922 752
905 736 913 752
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
830 579 859 603
840 587 848 603
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
841 498 866 522
849 506 857 522
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
839 416 868 440
849 424 857 440
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
888 920 917 944
898 928 906 944
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
893 1073 922 1097
903 1081 911 1097
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
897 1235 926 1259
907 1243 915 1259
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
973 304 1018 328
983 312 1007 328
3 Rbo
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
