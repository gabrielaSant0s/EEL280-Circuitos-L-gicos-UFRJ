CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.168350
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
99
13 Logic Switch~
5 246 1459 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3206 0 0
2
43729.7 0
0
13 Logic Switch~
5 195 1461 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 w
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9162 0 0
2
43729.7 1
0
13 Logic Switch~
5 145 1462 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9381 0 0
2
43729.7 2
0
13 Logic Switch~
5 89 1462 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 x
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4992 0 0
2
43729.7 3
0
13 Logic Switch~
5 290 85 0 1 11
0 92
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8456 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 226 83 0 1 11
0 75
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 W
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8342 0 0
2
5.89909e-315 5.26354e-315
0
13 Logic Switch~
5 174 82 0 1 11
0 77
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9685 0 0
2
5.89909e-315 5.30499e-315
0
13 Logic Switch~
5 116 82 0 1 11
0 80
0
0 0 21360 270
2 0V
-7 -21 7 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7318 0 0
2
5.89909e-315 5.32571e-315
0
8 2-In OR~
219 416 2878 0 3 22
0 15 14 12
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U27A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
3167 0 0
2
43729.9 0
0
9 2-In AND~
219 317 2928 0 3 22
0 18 23 20
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U40B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 42 0
1 U
3547 0 0
2
43729.9 5
0
9 2-In AND~
219 318 2975 0 3 22
0 22 21 19
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U40C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 42 0
1 U
9895 0 0
2
43729.9 4
0
8 2-In OR~
219 399 2948 0 3 22
0 20 19 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U39C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 41 0
1 U
5891 0 0
2
43729.9 1
0
8 3-In OR~
219 533 2878 0 4 22
0 11 12 13 17
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U38B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 40 0
1 U
8863 0 0
2
43729.9 0
0
8 2-In OR~
219 529 2692 0 3 22
0 30 29 24
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U39A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 41 0
1 U
393 0 0
2
43729.9 7
0
8 2-In OR~
219 444 2747 0 3 22
0 31 11 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 21 0
1 U
6476 0 0
2
43729.9 6
0
8 3-In OR~
219 437 2648 0 4 22
0 32 15 16 30
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U38A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 40 0
1 U
4421 0 0
2
43729.9 5
0
9 3-In AND~
219 356 2797 0 4 22
0 27 26 25 11
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U37A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 39 0
1 U
5341 0 0
2
43729.9 4
0
9 2-In AND~
219 358 2670 0 3 22
0 23 21 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U36B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 38 0
1 U
6395 0 0
2
43729.9 2
0
9 2-In AND~
219 358 2628 0 3 22
0 25 28 32
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U36A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 38 0
1 U
8741 0 0
2
43729.9 1
0
9 2-In AND~
219 357 2755 0 3 22
0 28 26 31
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U40D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 42 0
1 U
8261 0 0
2
43729.9 0
0
9 Inverter~
13 543 2501 0 2 22
0 4 33
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U34A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 36 0
1 U
7839 0 0
2
43729.9 5
0
9 2-In AND~
219 362 2574 0 3 22
0 23 22 16
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 35 0
1 U
8885 0 0
2
43729.9 4
0
9 4-In NOR~
219 459 2500 0 5 22
0 34 14 3 16 4
0
0 0 624 0
4 4002
-14 -24 14 -16
4 U35A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 37 0
1 U
3689 0 0
2
43729.9 2
0
9 2-In AND~
219 362 2459 0 3 22
0 23 26 34
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 35 0
1 U
3570 0 0
2
43729.9 1
0
9 2-In AND~
219 362 2497 0 3 22
0 22 28 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U23A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 25 0
1 U
9343 0 0
2
43729.9 0
0
9 2-In XOR~
219 322 2410 0 3 22
0 22 26 36
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U29C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 31 0
1 U
9817 0 0
2
43729.9 7
0
9 2-In AND~
219 417 2386 0 3 22
0 18 36 37
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U31A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 33 0
1 U
9129 0 0
2
43729.9 6
0
8 2-In OR~
219 497 2379 0 3 22
0 40 37 38
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U42B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 44 0
1 U
5573 0 0
2
43729.9 5
0
9 2-In AND~
219 414 2243 0 3 22
0 25 23 42
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U24A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
8151 0 0
2
43729.9 4
0
9 3-In AND~
219 415 2336 0 4 22
0 28 27 21 40
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U37C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 39 0
1 U
6375 0 0
2
43729.9 3
0
9 3-In AND~
219 414 2292 0 4 22
0 22 28 26 41
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U41B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 43 0
1 U
3122 0 0
2
43729.9 2
0
8 2-In OR~
219 482 2258 0 3 22
0 42 41 39
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U39D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 41 0
1 U
5719 0 0
2
43729.9 1
0
8 2-In OR~
219 575 2321 0 3 22
0 39 38 35
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U42A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 44 0
1 U
3569 0 0
2
43729.9 0
0
9 2-In AND~
219 301 2106 0 3 22
0 27 18 48
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U54D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 56 0
1 U
7688 0 0
2
43729.9 6
0
9 2-In AND~
219 300 2070 0 3 22
0 27 25 49
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U54B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 56 0
1 U
3316 0 0
2
43729.9 5
0
9 2-In AND~
219 302 2145 0 3 22
0 25 18 47
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U54C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 56 0
1 U
6741 0 0
2
43729.9 4
0
6 74136~
219 286 2197 0 3 22
0 23 26 46
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U55A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 57 0
1 U
593 0 0
2
43729.9 3
0
8 2-In OR~
219 358 2097 0 3 22
0 49 48 45
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U42C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 44 0
1 U
4132 0 0
2
43729.9 2
0
8 2-In OR~
219 359 2167 0 3 22
0 47 46 44
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U42D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 44 0
1 U
3574 0 0
2
43729.9 1
0
8 2-In OR~
219 432 2121 0 3 22
0 45 44 43
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U47A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 49 0
1 U
315 0 0
2
43729.9 0
0
6 74136~
219 290 2019 0 3 22
0 23 22 53
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U55B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 57 0
1 U
3889 0 0
2
43729.9 7
0
9 2-In AND~
219 365 2008 0 3 22
0 18 53 52
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U44A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 46 0
1 U
3545 0 0
2
43729.9 6
0
8 2-In OR~
219 587 1924 0 3 22
0 51 52 50
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U47D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 49 0
1 U
8315 0 0
2
43729.9 5
0
8 2-In OR~
219 496 1884 0 3 22
0 55 54 51
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U47C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 49 0
1 U
817 0 0
2
43729.9 4
0
9 2-In AND~
219 425 1923 0 3 22
0 28 56 54
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U50A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 52 0
1 U
9586 0 0
2
43729.9 3
0
9 2-In AND~
219 292 1970 0 3 22
0 25 27 57
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U25A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 27 0
1 U
3736 0 0
2
43729.9 2
0
8 2-In OR~
219 357 1949 0 3 22
0 21 57 56
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U47B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 49 0
1 U
4344 0 0
2
43729.9 1
0
9 2-In AND~
219 319 1894 0 3 22
0 27 21 55
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U49A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 51 0
1 U
5688 0 0
2
43729.9 0
0
8 3-In OR~
219 516 1668 0 4 22
0 62 61 60 66
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U46A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 48 0
1 U
7351 0 0
2
43729.8 0
0
8 2-In OR~
219 397 1575 0 3 22
0 65 64 62
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U45A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 47 0
1 U
392 0 0
2
43729.8 0
0
8 2-In OR~
219 400 1688 0 3 22
0 63 3 61
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U22A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
5788 0 0
2
43729.8 0
0
8 2-In OR~
219 394 1802 0 3 22
0 59 58 60
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U30D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
4290 0 0
2
43729.8 0
0
7 Ground~
168 950 2040 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3479 0 0
2
5.89909e-315 0
0
9 CC 7-Seg~
183 864 1875 0 17 19
10 66 50 43 35 33 24 17 105 2
1 0 0 0 1 1 1 2
0
0 0 21104 0
7 AMBERCC
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
886 0 0
2
5.89909e-315 0
0
7 Ground~
168 1422 1643 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8133 0 0
2
43729.7 25
0
4 LED~
171 1422 1611 0 2 2
10 67 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8564 0 0
2
43729.7 26
0
9 3-In AND~
219 320 1847 0 4 22
0 23 21 25 58
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 18 0
1 U
5876 0 0
2
43729.7 32
0
9 3-In AND~
219 321 1793 0 4 22
0 18 27 26 59
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 18 0
1 U
6693 0 0
2
43729.7 33
0
9 2-In AND~
219 324 1729 0 3 22
0 28 21 3
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 23 0
1 U
4551 0 0
2
43729.7 34
0
9 2-In AND~
219 324 1671 0 3 22
0 23 28 63
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5790 0 0
2
43729.7 35
0
9 2-In AND~
219 324 1615 0 3 22
0 26 22 64
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3845 0 0
2
43729.7 36
0
9 2-In AND~
219 322 1553 0 3 22
0 27 22 65
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8294 0 0
2
43729.7 37
0
9 Inverter~
13 175 1525 0 2 22
0 22 25
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U20A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 22 0
1 U
7344 0 0
2
43729.7 38
0
9 Inverter~
13 225 1526 0 2 22
0 18 28
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
3552 0 0
2
43729.7 39
0
9 Inverter~
13 59 1519 0 2 22
0 23 27
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
5966 0 0
2
43729.7 40
0
9 Inverter~
13 124 1520 0 2 22
0 26 21
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
3284 0 0
2
43729.7 41
0
7 Ground~
168 674 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
570 0 0
2
43729.7 42
0
9 CC 7-Seg~
183 607 384 0 17 19
10 74 73 72 71 70 69 68 106 2
1 1 1 1 1 1 0 2
0
0 0 21104 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3987 0 0
2
43729.7 43
0
8 2-In OR~
219 515 1013 0 3 22
0 80 82 85
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
7285 0 0
2
43729.7 44
0
8 2-In OR~
219 508 1124 0 3 22
0 84 83 81
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
3584 0 0
2
43729.7 45
0
8 2-In OR~
219 579 1073 0 3 22
0 85 81 68
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
3181 0 0
2
43729.7 46
0
9 2-In AND~
219 416 1034 0 3 22
0 75 76 82
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
3154 0 0
2
43729.7 47
0
9 2-In AND~
219 416 1092 0 3 22
0 77 78 84
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
3397 0 0
2
43729.7 48
0
9 2-In AND~
219 415 1151 0 3 22
0 75 79 83
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
3654 0 0
2
43729.7 49
0
8 2-In OR~
219 557 892 0 3 22
0 87 86 69
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
6959 0 0
2
43729.7 50
0
8 2-In OR~
219 482 930 0 3 22
0 89 88 86
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
3688 0 0
2
43729.7 51
0
8 2-In OR~
219 485 855 0 3 22
0 90 80 87
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
7228 0 0
2
43729.7 52
0
9 2-In AND~
219 409 832 0 3 22
0 77 79 90
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
6996 0 0
2
43729.7 53
0
9 2-In AND~
219 408 899 0 3 22
0 77 78 89
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
3550 0 0
2
43729.7 54
0
9 2-In AND~
219 405 958 0 3 22
0 78 79 88
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
9959 0 0
2
43729.7 55
0
9 2-In AND~
219 553 746 0 3 22
0 91 79 70
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
3122 0 0
2
43729.7 56
0
8 2-In OR~
219 446 717 0 3 22
0 76 75 91
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
5966 0 0
2
43729.7 57
0
9 3-In AND~
219 399 636 0 4 22
0 78 92 77 95
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 6 0
1 U
6493 0 0
2
5.89909e-315 5.34643e-315
0
8 3-In OR~
219 556 553 0 4 22
0 97 96 95 71
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
4738 0 0
2
5.89909e-315 5.3568e-315
0
8 3-In OR~
219 485 470 0 4 22
0 80 94 93 97
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
326 0 0
2
5.89909e-315 5.36716e-315
0
9 2-In AND~
219 403 481 0 3 22
0 79 75 94
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4484 0 0
2
5.89909e-315 5.37752e-315
0
9 2-In AND~
219 402 530 0 3 22
0 76 79 93
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
5360 0 0
2
5.89909e-315 5.38788e-315
0
9 2-In AND~
219 397 588 0 3 22
0 76 75 96
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
4548 0 0
2
5.89909e-315 5.39306e-315
0
8 2-In OR~
219 495 385 0 3 22
0 77 98 72
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
9370 0 0
2
5.89909e-315 5.39824e-315
0
8 2-In OR~
219 412 411 0 3 22
0 78 92 98
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3641 0 0
2
5.89909e-315 5.40342e-315
0
6 74266~
219 369 352 0 3 22
0 75 92 99
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7889 0 0
2
5.89909e-315 5.4086e-315
0
8 2-In OR~
219 491 303 0 3 22
0 76 99 73
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6725 0 0
2
5.89909e-315 5.41378e-315
0
8 2-In OR~
219 388 188 0 3 22
0 80 75 101
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3660 0 0
2
5.89909e-315 5.41896e-315
0
8 2-In OR~
219 485 221 0 3 22
0 101 100 74
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9613 0 0
2
5.89909e-315 5.42414e-315
0
6 74266~
219 390 264 0 3 22
0 77 92 100
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3418 0 0
2
5.89909e-315 5.42933e-315
0
9 Inverter~
13 260 136 0 2 22
0 92 79
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
3585 0 0
2
5.89909e-315 5.43192e-315
0
9 Inverter~
13 199 134 0 2 22
0 75 78
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
9150 0 0
2
5.89909e-315 5.43451e-315
0
9 Inverter~
13 143 131 0 2 22
0 77 76
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
367 0 0
2
5.89909e-315 5.4371e-315
0
9 Inverter~
13 82 132 0 2 22
0 80 102
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3420 0 0
2
5.89909e-315 5.43969e-315
0
210
3 0 3 0 0 8320 0 23 0 0 98 5
442 2505
391 2505
391 1834
352 1834
352 1729
5 1 4 0 0 8320 0 23 21 0 0 3
498 2500
498 2501
528 2501
1 0 11 0 0 16512 0 13 0 0 25 5
520 2869
470 2869
470 2837
421 2837
421 2756
3 2 12 0 0 4224 0 9 13 0 0 2
449 2878
521 2878
3 3 13 0 0 8320 0 12 13 0 0 4
432 2948
491 2948
491 2887
520 2887
2 0 14 0 0 8320 0 9 0 0 8 3
403 2887
387 2887
387 2496
1 0 15 0 0 4224 0 9 0 0 27 4
403 2869
403 2663
402 2663
402 2648
3 2 14 0 0 0 0 25 23 0 0 4
383 2497
387 2497
387 2496
442 2496
3 0 16 0 0 8320 0 16 0 0 36 3
424 2657
409 2657
409 2574
7 4 17 0 0 4224 0 54 13 0 0 3
879 1911
879 2878
566 2878
1 0 18 0 0 4096 0 10 0 0 129 2
293 2919
246 2919
3 2 19 0 0 4224 0 11 12 0 0 4
339 2975
367 2975
367 2957
386 2957
3 1 20 0 0 4224 0 10 12 0 0 4
338 2928
366 2928
366 2939
386 2939
2 0 21 0 0 4096 0 11 0 0 122 2
294 2984
127 2984
1 0 22 0 0 4096 0 11 0 0 130 2
294 2966
195 2966
2 0 23 0 0 4096 0 10 0 0 132 2
293 2937
89 2937
6 3 24 0 0 4224 0 54 14 0 0 3
873 1911
873 2692
562 2692
3 0 25 0 0 4096 0 17 0 0 123 2
332 2806
178 2806
2 0 26 0 0 4096 0 17 0 0 131 2
332 2797
145 2797
1 0 27 0 0 4096 0 17 0 0 121 2
332 2788
62 2788
2 0 26 0 0 4096 0 20 0 0 131 2
333 2764
145 2764
1 0 28 0 0 4096 0 20 0 0 124 2
333 2746
228 2746
3 2 29 0 0 8320 0 15 14 0 0 4
477 2747
488 2747
488 2701
516 2701
4 1 30 0 0 8320 0 16 14 0 0 4
470 2648
487 2648
487 2683
516 2683
4 2 11 0 0 0 0 17 15 0 0 4
377 2797
415 2797
415 2756
431 2756
3 1 31 0 0 8320 0 20 15 0 0 3
378 2755
378 2738
431 2738
3 2 15 0 0 0 0 18 16 0 0 4
379 2670
397 2670
397 2648
425 2648
3 1 32 0 0 12416 0 19 16 0 0 4
379 2628
398 2628
398 2639
424 2639
2 0 21 0 0 4096 0 18 0 0 122 2
334 2679
127 2679
1 0 23 0 0 4096 0 18 0 0 132 2
334 2661
89 2661
2 0 28 0 0 4096 0 19 0 0 124 2
334 2637
228 2637
1 0 25 0 0 4096 0 19 0 0 123 2
334 2619
178 2619
5 2 33 0 0 4224 0 54 21 0 0 3
867 1911
867 2501
564 2501
2 0 28 0 0 4096 0 25 0 0 124 2
338 2506
228 2506
1 0 22 0 0 4096 0 25 0 0 130 2
338 2488
195 2488
3 4 16 0 0 0 0 22 23 0 0 4
383 2574
435 2574
435 2514
442 2514
3 1 34 0 0 12416 0 24 23 0 0 4
383 2459
412 2459
412 2487
442 2487
2 0 22 0 0 0 0 22 0 0 130 2
338 2583
195 2583
1 0 23 0 0 4096 0 22 0 0 132 2
338 2565
89 2565
2 0 26 0 0 4096 0 24 0 0 131 2
338 2468
145 2468
1 0 23 0 0 0 0 24 0 0 132 2
338 2450
89 2450
4 3 35 0 0 4224 0 54 33 0 0 3
861 1911
861 2321
608 2321
3 2 36 0 0 12416 0 26 27 0 0 4
355 2410
372 2410
372 2395
393 2395
2 0 26 0 0 0 0 26 0 0 131 2
306 2419
145 2419
1 0 22 0 0 0 0 26 0 0 130 2
306 2401
195 2401
1 0 18 0 0 4096 0 27 0 0 129 2
393 2377
246 2377
3 2 37 0 0 4224 0 27 28 0 0 4
438 2386
476 2386
476 2388
484 2388
3 2 38 0 0 8320 0 28 33 0 0 4
530 2379
535 2379
535 2330
562 2330
3 1 39 0 0 8320 0 32 33 0 0 4
515 2258
535 2258
535 2312
562 2312
4 1 40 0 0 8320 0 30 28 0 0 4
436 2336
452 2336
452 2370
484 2370
4 2 41 0 0 8320 0 31 32 0 0 4
435 2292
452 2292
452 2267
469 2267
3 1 42 0 0 12416 0 29 32 0 0 4
435 2243
448 2243
448 2249
469 2249
3 0 21 0 0 4096 0 30 0 0 122 2
391 2345
127 2345
2 0 27 0 0 4096 0 30 0 0 121 2
391 2336
62 2336
1 0 28 0 0 4096 0 30 0 0 124 2
391 2327
228 2327
3 0 26 0 0 4096 0 31 0 0 131 2
390 2301
145 2301
2 0 28 0 0 0 0 31 0 0 124 2
390 2292
228 2292
1 0 22 0 0 4096 0 31 0 0 130 2
390 2283
195 2283
2 0 23 0 0 4096 0 29 0 0 132 2
390 2252
89 2252
1 0 25 0 0 4096 0 29 0 0 123 2
390 2234
178 2234
3 3 43 0 0 8320 0 54 40 0 0 3
855 1911
855 2121
465 2121
2 0 26 0 0 0 0 37 0 0 131 2
270 2206
145 2206
1 0 23 0 0 0 0 37 0 0 132 2
270 2188
89 2188
2 0 18 0 0 0 0 36 0 0 129 2
278 2154
246 2154
1 0 25 0 0 0 0 36 0 0 123 2
278 2136
178 2136
2 0 18 0 0 0 0 34 0 0 129 2
277 2115
246 2115
1 0 27 0 0 0 0 34 0 0 121 2
277 2097
62 2097
2 0 25 0 0 0 0 35 0 0 123 2
276 2079
178 2079
1 0 27 0 0 0 0 35 0 0 121 2
276 2061
62 2061
3 2 44 0 0 8320 0 39 40 0 0 4
392 2167
402 2167
402 2130
419 2130
3 1 45 0 0 12416 0 38 40 0 0 4
391 2097
403 2097
403 2112
419 2112
3 2 46 0 0 8320 0 37 39 0 0 4
319 2197
336 2197
336 2176
346 2176
3 1 47 0 0 4224 0 36 39 0 0 4
323 2145
336 2145
336 2158
346 2158
3 2 48 0 0 4224 0 34 38 0 0 2
322 2106
345 2106
3 1 49 0 0 8320 0 35 38 0 0 4
321 2070
333 2070
333 2088
345 2088
2 3 50 0 0 8320 0 54 43 0 0 3
849 1911
849 1924
620 1924
3 1 51 0 0 8320 0 44 43 0 0 4
529 1884
546 1884
546 1915
574 1915
3 2 52 0 0 12416 0 42 43 0 0 4
386 2008
475 2008
475 1933
574 1933
3 2 53 0 0 8320 0 41 42 0 0 3
323 2019
323 2017
341 2017
1 0 18 0 0 0 0 42 0 0 129 2
341 1999
246 1999
2 0 22 0 0 0 0 41 0 0 130 2
274 2028
195 2028
1 0 23 0 0 0 0 41 0 0 132 2
274 2010
89 2010
3 2 54 0 0 8320 0 45 44 0 0 4
446 1923
467 1923
467 1893
483 1893
3 1 55 0 0 4224 0 48 44 0 0 4
340 1894
455 1894
455 1875
483 1875
3 2 56 0 0 8320 0 47 45 0 0 3
390 1949
401 1949
401 1932
1 0 28 0 0 4096 0 45 0 0 124 2
401 1914
228 1914
3 2 57 0 0 12416 0 46 47 0 0 4
313 1970
325 1970
325 1958
344 1958
1 0 21 0 0 0 0 47 0 0 122 2
344 1940
127 1940
2 0 27 0 0 0 0 46 0 0 121 2
268 1979
62 1979
1 0 25 0 0 0 0 46 0 0 123 2
268 1961
178 1961
2 0 21 0 0 0 0 48 0 0 122 2
295 1903
127 1903
1 0 27 0 0 0 0 48 0 0 121 2
295 1885
62 1885
4 2 58 0 0 4224 0 57 52 0 0 4
341 1847
377 1847
377 1811
381 1811
4 1 59 0 0 4224 0 58 52 0 0 2
342 1793
381 1793
3 3 60 0 0 8320 0 52 49 0 0 4
427 1802
494 1802
494 1677
503 1677
3 2 61 0 0 4224 0 51 49 0 0 4
433 1688
483 1688
483 1668
504 1668
3 1 62 0 0 8320 0 50 49 0 0 4
430 1575
465 1575
465 1659
503 1659
3 2 3 0 0 128 0 59 51 0 0 4
345 1729
379 1729
379 1697
387 1697
3 1 63 0 0 4224 0 60 51 0 0 4
345 1671
379 1671
379 1679
387 1679
3 2 64 0 0 4224 0 61 50 0 0 4
345 1615
376 1615
376 1584
384 1584
3 1 65 0 0 12416 0 62 50 0 0 4
343 1553
357 1553
357 1566
384 1566
4 0 66 0 0 12288 0 49 0 0 104 4
549 1668
581 1668
581 1711
654 1711
9 1 2 0 0 8320 0 54 53 0 0 3
864 1833
950 1833
950 2034
0 1 66 0 0 8320 0 0 54 0 0 5
651 1711
758 1711
758 1921
843 1921
843 1911
3 1 67 0 0 4224 0 0 56 0 0 3
1385 1572
1422 1572
1422 1601
1 2 2 0 0 0 0 55 56 0 0 2
1422 1637
1422 1621
3 0 25 0 0 0 0 57 0 0 123 2
296 1856
178 1856
2 0 21 0 0 0 0 57 0 0 122 2
296 1847
127 1847
1 0 23 0 0 0 0 60 0 0 132 2
300 1662
89 1662
1 0 23 0 0 0 0 57 0 0 132 2
296 1838
89 1838
3 0 26 0 0 0 0 58 0 0 131 2
297 1802
145 1802
2 0 27 0 0 0 0 58 0 0 121 2
297 1793
62 1793
1 0 18 0 0 0 0 58 0 0 129 2
297 1784
246 1784
2 0 21 0 0 0 0 59 0 0 122 2
300 1738
127 1738
1 0 28 0 0 0 0 59 0 0 124 2
300 1720
228 1720
2 0 28 0 0 0 0 60 0 0 124 2
300 1680
228 1680
2 0 22 0 0 0 0 61 0 0 130 2
300 1624
195 1624
1 0 26 0 0 0 0 61 0 0 131 2
300 1606
145 1606
2 0 22 0 0 0 0 62 0 0 130 2
298 1562
195 1562
0 1 27 0 0 0 0 0 62 121 0 3
62 1543
62 1544
298 1544
2 0 27 0 0 4224 0 65 0 0 0 2
62 1537
62 3263
2 0 21 0 0 4224 0 66 0 0 0 2
127 1538
127 3262
2 0 25 0 0 4224 0 63 0 0 0 2
178 1543
178 3263
2 0 28 0 0 4224 0 64 0 0 0 2
228 1544
228 3264
1 0 18 0 0 0 0 64 0 0 129 3
228 1508
228 1483
246 1483
1 0 22 0 0 0 0 63 0 0 130 3
178 1507
178 1483
195 1483
1 0 26 0 0 0 0 66 0 0 131 3
127 1502
127 1484
145 1484
1 0 23 0 0 0 0 65 0 0 132 3
62 1501
62 1486
89 1486
1 0 18 0 0 4224 0 1 0 0 0 2
246 1471
246 3265
1 0 22 0 0 4224 0 2 0 0 0 2
195 1473
195 3264
1 0 26 0 0 4224 0 3 0 0 0 2
145 1474
145 3264
1 0 23 0 0 4224 0 4 0 0 0 2
89 1474
89 3264
7 3 68 0 0 4224 0 68 71 0 0 3
622 420
622 1073
612 1073
6 3 69 0 0 4224 0 68 75 0 0 3
616 420
616 892
590 892
5 3 70 0 0 4224 0 68 81 0 0 3
610 420
610 746
574 746
4 4 71 0 0 4224 0 68 84 0 0 3
604 420
604 553
589 553
3 3 72 0 0 8320 0 68 89 0 0 5
598 420
598 430
541 430
541 385
528 385
2 3 73 0 0 12416 0 68 92 0 0 5
592 420
592 425
537 425
537 303
524 303
1 3 74 0 0 8320 0 68 94 0 0 4
586 420
533 420
533 221
518 221
1 9 2 0 0 0 0 67 68 0 0 4
674 426
674 330
607 330
607 342
1 0 75 0 0 4096 0 72 0 0 203 2
392 1025
226 1025
2 0 76 0 0 4096 0 72 0 0 206 2
392 1043
146 1043
1 0 77 0 0 4096 0 73 0 0 207 2
392 1083
174 1083
2 0 78 0 0 4096 0 73 0 0 202 2
392 1101
202 1101
2 0 79 0 0 4096 0 74 0 0 200 2
391 1160
263 1160
1 0 75 0 0 0 0 74 0 0 203 2
391 1142
226 1142
1 0 80 0 0 4096 0 69 0 0 210 2
502 1004
116 1004
3 2 81 0 0 8320 0 70 71 0 0 4
541 1124
558 1124
558 1082
566 1082
3 2 82 0 0 4224 0 72 69 0 0 4
437 1034
471 1034
471 1022
502 1022
3 2 83 0 0 4224 0 74 70 0 0 4
436 1151
476 1151
476 1133
495 1133
3 1 84 0 0 4224 0 73 70 0 0 4
437 1092
476 1092
476 1115
495 1115
3 1 85 0 0 4224 0 69 71 0 0 3
548 1013
548 1064
566 1064
2 0 79 0 0 0 0 80 0 0 200 2
381 967
263 967
2 0 78 0 0 0 0 79 0 0 202 2
384 908
202 908
1 0 78 0 0 0 0 80 0 0 202 2
381 949
202 949
2 0 79 0 0 0 0 78 0 0 200 2
385 841
263 841
1 0 77 0 0 0 0 78 0 0 207 2
385 823
174 823
2 0 80 0 0 0 0 77 0 0 210 2
472 864
116 864
3 2 86 0 0 8320 0 76 75 0 0 4
515 930
536 930
536 901
544 901
3 1 87 0 0 8320 0 77 75 0 0 4
518 855
536 855
536 883
544 883
3 2 88 0 0 4224 0 80 76 0 0 4
426 958
461 958
461 939
469 939
3 1 89 0 0 4224 0 79 76 0 0 4
429 899
461 899
461 921
469 921
3 1 90 0 0 8320 0 78 77 0 0 3
430 832
430 846
472 846
0 1 77 0 0 0 0 0 79 207 0 2
174 890
384 890
0 2 79 0 0 4096 0 0 81 200 0 4
263 781
513 781
513 755
529 755
3 1 91 0 0 4224 0 82 81 0 0 4
479 717
512 717
512 737
529 737
0 2 75 0 0 4096 0 0 82 203 0 4
226 741
396 741
396 726
433 726
0 1 76 0 0 4096 0 0 82 206 0 4
146 693
396 693
396 708
433 708
3 0 77 0 0 0 0 83 0 0 207 2
375 645
174 645
2 0 92 0 0 4096 0 83 0 0 199 2
375 636
290 636
1 0 78 0 0 0 0 83 0 0 202 2
375 627
202 627
2 0 75 0 0 0 0 88 0 0 203 2
373 597
226 597
1 0 76 0 0 0 0 88 0 0 206 2
373 579
146 579
2 0 79 0 0 0 0 87 0 0 200 2
378 539
263 539
1 0 79 0 0 0 0 86 0 0 200 2
379 472
263 472
1 0 76 0 0 0 0 87 0 0 206 2
378 521
146 521
2 0 75 0 0 0 0 86 0 0 203 2
379 490
226 490
3 3 93 0 0 8320 0 87 85 0 0 4
423 530
452 530
452 479
472 479
3 2 94 0 0 12416 0 86 85 0 0 4
424 481
440 481
440 470
473 470
1 0 80 0 0 0 0 85 0 0 210 2
472 461
116 461
4 3 95 0 0 4224 0 83 84 0 0 4
420 636
520 636
520 562
543 562
3 2 96 0 0 4224 0 88 84 0 0 4
418 588
495 588
495 553
544 553
4 1 97 0 0 8320 0 85 84 0 0 4
518 470
535 470
535 544
543 544
1 0 78 0 0 4096 0 90 0 0 202 2
399 402
202 402
2 0 92 0 0 4096 0 90 0 0 199 2
399 420
290 420
1 0 77 0 0 4096 0 89 0 0 207 2
482 376
174 376
3 2 98 0 0 4224 0 90 89 0 0 4
445 411
474 411
474 394
482 394
2 0 92 0 0 0 0 91 0 0 199 2
353 361
290 361
1 0 75 0 0 0 0 91 0 0 203 2
353 343
226 343
1 0 76 0 0 4096 0 92 0 0 206 2
478 294
146 294
3 2 99 0 0 8320 0 91 92 0 0 3
408 352
408 312
478 312
2 0 92 0 0 0 0 95 0 0 199 2
374 273
290 273
1 0 80 0 0 0 0 93 0 0 210 2
375 179
116 179
3 2 100 0 0 4224 0 95 94 0 0 4
429 264
464 264
464 230
472 230
0 1 77 0 0 0 0 0 95 207 0 4
174 220
367 220
367 255
374 255
0 2 75 0 0 0 0 0 93 203 0 4
226 260
349 260
349 197
375 197
3 1 101 0 0 4224 0 93 94 0 0 4
421 188
452 188
452 212
472 212
0 1 92 0 0 0 0 0 96 199 0 3
290 109
263 109
263 118
1 0 92 0 0 4224 0 5 0 0 0 2
290 97
290 1209
2 0 79 0 0 4224 0 96 0 0 0 2
263 154
263 1212
1 0 75 0 0 0 0 97 0 0 203 2
202 116
226 116
2 0 78 0 0 4224 0 97 0 0 0 2
202 152
202 1215
1 0 75 0 0 4224 0 6 0 0 0 2
226 95
226 1212
1 0 77 0 0 0 0 98 0 0 207 2
146 113
174 113
1 0 80 0 0 0 0 99 0 0 210 2
85 114
116 114
2 0 76 0 0 4224 0 98 0 0 0 2
146 149
146 1215
1 0 77 0 0 4224 0 7 0 0 0 2
174 94
174 1214
1 0 77 0 0 0 0 7 0 0 0 2
174 94
174 656
2 0 102 0 0 4224 0 99 0 0 0 2
85 150
85 1217
1 0 80 0 0 4224 0 8 0 0 0 2
116 94
116 1216
18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
565 2837 590 2861
573 2845 581 2861
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
567 2655 592 2679
575 2663 583 2679
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
563 2471 588 2495
571 2479 579 2495
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
614 2285 639 2309
622 2293 630 2309
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
485 2076 510 2100
493 2084 501 2100
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
348 2112 377 2136
358 2120 366 2136
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
612 1875 637 1899
620 1883 628 1899
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 37
245 1377 562 1401
255 1385 551 1401
37 Decodificador hexadecimal 7 segmentos
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
239 11 492 35
249 19 481 35
29 Decodificador BCD 7 segmentos
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 5 55 29
28 13 44 29
2 a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
654 1669 683 1693
664 1677 672 1693
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 1006 614 1030
595 1014 603 1030
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
581 844 610 868
591 852 599 868
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
576 691 605 715
586 699 594 715
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
527 187 556 211
537 195 545 211
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
529 269 554 293
537 277 545 293
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
518 350 547 374
528 358 536 374
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 499 610 523
593 507 601 523
1 d
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
