CircuitMaker Text
5.6
Probes: 1
A_1
Operating Point
0 273 233 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
360 670 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
1083179026 0
0
6 Title:
5 Name:
0
0
0
39
13 Logic Switch~
5 852 943 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43723 0
0
13 Logic Switch~
5 855 987 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43723 1
0
13 Logic Switch~
5 858 767 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43723 2
0
13 Logic Switch~
5 859 723 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43723 3
0
13 Logic Switch~
5 877 507 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
43723 4
0
13 Logic Switch~
5 878 463 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
43723 5
0
13 Logic Switch~
5 903 210 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
43723 6
0
13 Logic Switch~
5 902 254 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
43723 7
0
13 Logic Switch~
5 246 747 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
43723 8
0
13 Logic Switch~
5 248 503 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
43723 9
0
13 Logic Switch~
5 247 547 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
43723 10
0
13 Logic Switch~
5 250 275 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
43723 11
0
13 Logic Switch~
5 251 231 0 1 11
0 27
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
43723 12
0
5 4030~
219 1004 961 0 3 22
0 11 10 12
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
4597 0 0
2
43723 13
0
7 Ground~
168 1138 1028 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
43723 14
0
4 LED~
171 1137 977 0 2 2
10 9 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3670 0 0
2
43723 15
0
10 2-In XNOR~
219 1003 741 0 3 22
0 14 13 15
0
0 0 608 0
4 4077
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
5616 0 0
2
43723 16
0
4 LED~
171 1140 757 0 2 2
10 8 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9323 0 0
2
43723 17
0
7 Ground~
168 1141 808 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
43723 18
0
10 2-In NAND~
219 1007 480 0 3 22
0 18 17 16
0
0 0 608 0
5 74F37
-10 -24 25 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3108 0 0
2
43723 19
0
4 LED~
171 1159 497 0 2 2
10 7 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4299 0 0
2
43723 20
0
7 Ground~
168 1160 548 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
43723 21
0
5 4001~
219 1020 227 0 3 22
0 20 19 21
0
0 0 608 0
4 4001
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 4 0
1 U
7876 0 0
2
43723 22
0
7 Ground~
168 1185 295 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
43723 23
0
4 LED~
171 1184 244 0 2 2
10 5 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9172 0 0
2
43723 24
0
9 Inverter~
13 377 764 0 2 22
0 22 3
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
7100 0 0
2
43723 25
0
4 LED~
171 527 781 0 2 2
10 3 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3820 0 0
2
43723 26
0
7 Ground~
168 528 832 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7678 0 0
2
43723 27
0
9 2-In AND~
219 378 520 0 3 22
0 25 24 23
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
961 0 0
2
43723 28
0
7 Ground~
168 530 588 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
43723 29
0
4 LED~
171 529 537 0 2 2
10 6 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3409 0 0
2
43723 30
0
8 2-In OR~
219 372 248 0 3 22
0 27 26 4
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3951 0 0
2
5.89908e-315 0
0
4 LED~
171 532 265 0 2 2
10 4 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8885 0 0
2
43723 31
0
7 Ground~
168 533 316 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3780 0 0
2
43723 32
0
9 Resistor~
219 460 519 0 2 5
0 23 6
0
0 0 864 0
3 200
-11 -14 10 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
5.89908e-315 0
0
9 Resistor~
219 1121 227 0 2 5
0 21 5
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9442 0 0
2
43723 33
0
9 Resistor~
219 1085 480 0 2 5
0 16 7
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9424 0 0
2
43723 34
0
9 Resistor~
219 1089 740 0 2 5
0 15 8
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
43723 35
0
9 Resistor~
219 1094 960 0 2 5
0 12 9
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
43723 36
0
36
2 1 3 0 0 4224 0 26 27 0 0 3
398 764
527 764
527 771
3 1 4 0 0 4224 0 32 33 0 0 3
405 248
532 248
532 255
2 1 5 0 0 4224 0 36 25 0 0 3
1139 227
1184 227
1184 234
2 1 6 0 0 8320 0 35 31 0 0 4
478 519
478 520
529 520
529 527
2 1 7 0 0 4224 0 37 21 0 0 3
1103 480
1159 480
1159 487
2 1 8 0 0 4224 0 38 18 0 0 3
1107 740
1140 740
1140 747
2 1 9 0 0 4224 0 39 16 0 0 3
1112 960
1137 960
1137 967
1 2 10 0 0 4224 0 2 14 0 0 4
867 987
980 987
980 970
988 970
1 1 11 0 0 4224 0 1 14 0 0 4
864 943
980 943
980 952
988 952
3 1 12 0 0 12416 0 14 39 0 0 4
1037 961
1039 961
1039 960
1076 960
1 2 2 0 0 8320 0 15 16 0 0 3
1138 1022
1137 1022
1137 987
2 0 13 0 0 4096 0 17 0 0 16 2
987 750
960 750
1 0 14 0 0 4096 0 17 0 0 17 3
987 732
961 731
960 731
3 1 15 0 0 8320 0 17 38 0 0 3
1042 741
1042 740
1071 740
1 2 2 0 0 0 0 19 18 0 0 3
1141 802
1140 802
1140 767
1 0 13 0 0 4224 0 3 0 0 0 4
870 767
960 767
960 749
966 749
1 0 14 0 0 4224 0 4 0 0 0 4
871 723
960 723
960 731
966 731
3 1 16 0 0 4224 0 20 37 0 0 2
1034 480
1067 480
1 2 2 0 0 0 0 22 21 0 0 3
1160 542
1159 542
1159 507
1 2 17 0 0 4224 0 5 20 0 0 4
889 507
979 507
979 489
983 489
1 1 18 0 0 4224 0 6 20 0 0 4
890 463
979 463
979 471
983 471
2 0 19 0 0 0 0 23 0 0 26 2
1007 236
1007 236
1 0 20 0 0 0 0 23 0 0 27 2
1007 218
1007 218
3 1 21 0 0 4224 0 23 36 0 0 2
1059 227
1103 227
1 2 2 0 0 0 0 24 25 0 0 3
1185 289
1184 289
1184 254
1 0 19 0 0 4224 0 8 0 0 0 4
914 254
1004 254
1004 236
1011 236
1 0 20 0 0 4224 0 7 0 0 0 4
915 210
1004 210
1004 218
1011 218
1 1 22 0 0 4224 0 9 26 0 0 4
258 747
354 747
354 764
362 764
1 2 2 0 0 0 0 28 27 0 0 3
528 826
527 826
527 791
3 1 23 0 0 4224 0 29 35 0 0 3
399 520
442 520
442 519
1 2 2 0 0 0 0 30 31 0 0 3
530 582
529 582
529 547
1 2 24 0 0 4224 0 11 29 0 0 4
259 547
349 547
349 529
354 529
1 1 25 0 0 4224 0 10 29 0 0 4
260 503
349 503
349 511
354 511
1 2 2 0 0 0 0 34 33 0 0 3
533 310
532 310
532 275
1 2 26 0 0 4224 0 12 32 0 0 4
262 275
352 275
352 257
359 257
1 1 27 0 0 4224 0 13 32 0 0 4
263 231
352 231
352 239
359 239
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 79
1234 902 1375 1066
1244 910 1364 1038
79 
     XOR 

A B | A'B + AB' 
0 0 | 	  0
0 1 | 	  1
1 0 | 	  1
1 1 | 	  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 80
1237 682 1378 846
1247 690 1367 818
80 
     XNOR 

A B | (AB)'+ AB 
0 0 | 	  1
0 1 | 	  0
1 0 | 	  0
1 1 | 	  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 68
1281 169 1414 333
1291 177 1403 305
68 
   NOR 

A B | (A + B)' 
0 0 | 	1
0 1 | 	0
1 0 | 	0
1 1 | 	0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
982 91 1155 115
992 99 1144 115
19 FUNCOES SECUNDARIAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
412 82 569 106
422 90 558 106
17 FUNCOES PRIMARIAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
631 659 716 803
641 667 705 779
40 
   NOT 

A  |  A' 
0  |  0
1  |  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 64
636 143 745 307
646 151 734 279
64 
   OR 

A B | A + B 
0 0 | 	0
0 1 | 	1
1 0 | 	1
1 1 | 	1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 65
623 455 732 619
633 463 721 591
65 
   AND 

A B | A . B 
0 0 | 	0
0 1 | 	0
1 0 | 	0
1 1 | 	1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 68
1256 422 1389 586
1266 430 1378 558
68 
   NAND

A B | (A . B)' 
0 0 | 	1
0 1 | 	1
1 0 | 	1
1 1 | 	0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
