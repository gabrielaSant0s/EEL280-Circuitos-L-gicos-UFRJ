CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 27 153 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-1 -13 13 -5
1 D
-13 -16 -6 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43739 0
0
13 Logic Switch~
5 29 124 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43739 1
0
13 Logic Switch~
5 28 88 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
43739 2
0
13 Logic Switch~
5 30 56 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43739 3
0
5 4073~
219 293 304 0 4 22
0 4 2 3 17
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 5 0
1 U
8157 0 0
2
5.8991e-315 0
0
14 Logic Display~
6 645 231 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
43739 4
0
14 Logic Display~
6 679 231 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -19 7 -11
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
43739 5
0
14 Logic Display~
6 712 231 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
43739 6
0
14 Logic Display~
6 741 231 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
43739 7
0
5 4081~
219 545 474 0 3 22
0 8 5 19
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
972 0 0
2
43739 8
0
5 4049~
219 100 236 0 2 22
0 5 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-1 -13 20 -5
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
3472 0 0
2
43739 9
0
5 4049~
219 101 216 0 2 22
0 3 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
3 -12 24 -4
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
9998 0 0
2
43739 10
0
8 4-In OR~
219 551 414 0 5 22
0 11 6 10 9 7
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
3536 0 0
2
43739 11
0
5 4073~
219 273 379 0 4 22
0 14 8 3 11
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 5 0
1 U
4597 0 0
2
43739 12
0
5 4073~
219 219 449 0 4 22
0 4 2 5 10
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U5A
9 -19 30 -11
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
3835 0 0
2
43739 13
0
5 4073~
219 272 347 0 4 22
0 4 3 13 16
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2C
8 -20 29 -12
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
3670 0 0
2
43739 14
0
5 4071~
219 440 332 0 3 22
0 17 16 15
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
5616 0 0
2
43739 15
0
5 4049~
219 101 196 0 2 22
0 8 2
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
0 -14 21 -6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
9323 0 0
2
43739 16
0
5 4073~
219 233 410 0 4 22
0 8 3 13 6
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
8 -23 29 -15
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
317 0 0
2
43739 17
0
5 4049~
219 101 176 0 2 22
0 4 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
1 -14 22 -6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3108 0 0
2
43739 18
0
5 4073~
219 220 482 0 4 22
0 4 12 5 9
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
7 -17 28 -9
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
4299 0 0
2
43739 19
0
5 4082~
219 227 261 0 5 22
0 4 8 3 5 18
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
9672 0 0
2
43739 20
0
47
0 2 2 0 0 4096 0 0 15 38 0 3
155 196
155 449
195 449
3 0 3 0 0 4096 0 14 0 0 3 2
249 388
67 388
0 0 3 0 0 0 0 0 0 27 20 2
67 345
67 410
2 0 2 0 0 0 0 5 0 0 38 3
269 304
256 304
256 196
1 0 4 0 0 4096 0 5 0 0 28 2
269 295
49 295
0 2 5 0 0 4096 0 0 10 44 0 3
353 153
353 483
521 483
2 4 6 0 0 4224 0 13 19 0 0 2
534 410
254 410
5 1 7 0 0 8320 0 13 8 0 0 3
584 414
712 414
712 249
1 0 8 0 0 8192 0 10 0 0 46 3
521 465
372 465
372 88
4 4 9 0 0 4224 0 13 21 0 0 4
534 428
288 428
288 482
241 482
4 3 10 0 0 12416 0 15 13 0 0 4
240 449
271 449
271 419
534 419
4 1 11 0 0 4224 0 14 13 0 0 4
294 379
485 379
485 401
534 401
3 0 5 0 0 0 0 21 0 0 16 3
196 491
74 491
74 458
0 2 12 0 0 4096 0 0 21 37 0 3
185 216
185 482
196 482
0 1 4 0 0 0 0 0 21 18 0 3
49 440
49 473
196 473
3 0 5 0 0 0 0 15 0 0 40 3
195 458
74 458
74 234
0 1 8 0 0 0 0 0 19 21 0 3
58 397
58 401
209 401
0 1 4 0 0 0 0 0 15 28 0 3
49 339
49 440
195 440
0 3 13 0 0 8192 0 0 19 26 0 3
126 357
126 419
209 419
2 0 3 0 0 0 0 19 0 0 0 3
209 410
67 410
67 407
0 2 8 0 0 0 0 0 14 42 0 5
58 196
58 397
58 397
58 379
249 379
0 1 14 0 0 4096 0 0 14 39 0 3
142 176
142 370
249 370
3 1 15 0 0 4224 0 17 7 0 0 3
473 332
679 332
679 249
4 2 16 0 0 12416 0 16 17 0 0 4
293 347
343 347
343 341
427 341
4 1 17 0 0 12416 0 5 17 0 0 4
314 304
342 304
342 323
427 323
0 3 13 0 0 16400 0 0 16 36 0 5
126 236
126 357
126 357
126 356
248 356
0 2 3 0 0 0 0 0 16 29 0 3
67 322
67 347
248 347
0 1 4 0 0 0 0 0 16 43 0 5
49 176
49 339
49 339
49 338
248 338
3 0 3 0 0 4096 0 5 0 0 41 5
269 313
67 313
67 322
65 322
65 216
5 1 18 0 0 4224 0 22 6 0 0 3
248 261
645 261
645 249
3 1 19 0 0 8320 0 10 9 0 0 3
566 474
741 474
741 249
4 0 5 0 0 0 0 22 0 0 44 3
203 275
176 275
176 153
3 0 3 0 0 0 0 22 0 0 45 3
203 266
163 266
163 124
2 0 8 0 0 0 0 22 0 0 46 3
203 257
150 257
150 88
1 0 4 0 0 0 0 22 0 0 47 3
203 248
136 248
136 56
2 0 13 0 0 4224 0 11 0 0 0 2
121 236
608 236
2 0 12 0 0 4224 0 12 0 0 0 2
122 216
608 216
2 0 2 0 0 4224 0 18 0 0 0 2
122 196
608 196
2 0 14 0 0 4224 0 20 0 0 0 2
122 176
608 176
0 1 5 0 0 0 0 0 11 44 0 3
74 153
74 236
85 236
1 0 3 0 0 0 0 12 0 0 45 3
86 216
64 216
64 124
1 0 8 0 0 0 0 18 0 0 46 3
86 196
57 196
57 88
1 0 4 0 0 0 0 20 0 0 47 3
86 176
48 176
48 56
1 0 5 0 0 4224 0 1 0 0 0 2
39 153
608 153
1 0 3 0 0 4224 0 2 0 0 0 2
41 124
608 124
1 0 8 0 0 4224 0 3 0 0 0 2
40 88
610 88
1 0 4 0 0 4224 0 4 0 0 0 2
42 56
610 56
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
