CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 110 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.253589 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
154
13 Logic Switch~
5 300 829 0 1 11
0 129
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 UD
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8856 0 0
2
43796 0
0
14 Logic Display~
6 496 199 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
469 0 0
2
43796 0
0
14 Logic Display~
6 275 207 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4529 0 0
2
5.89917e-315 0
0
2 +V
167 1350 852 0 1 3
0 14
0
0 0 54256 180
2 5V
-12 7 2 15
2 V5
-21 -10 -7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
88 0 0
2
43796 1
0
7 Ground~
168 1374 852 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3894 0 0
2
43796 2
0
6 74LS85
106 1510 794 0 14 29
0 10 11 12 13 2 2 2 14 140
141 142 5 6 7
0
0 0 5104 0
5 74F85
-18 -52 17 -44
3 U15
-11 -62 10 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6890 0 0
2
43796 3
0
6 74LS85
106 1510 688 0 14 29
0 2 2 8 9 2 2 14 2 5
6 7 143 4 3
0
0 0 5104 0
5 74F85
-18 -52 17 -44
3 U13
-11 -62 10 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3257 0 0
2
43796 4
0
7 Ground~
168 160 1301 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6612 0 0
2
43796 5
0
12 Hex Display~
7 75 1299 0 18 19
10 26 29 25 2 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP7
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3556 0 0
2
43796 6
0
8 2-In OR~
219 202 1455 0 3 22
0 28 27 26
0
0 0 624 512
5 74F32
-18 -24 17 -16
4 U11A
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
9143 0 0
2
43796 7
0
9 2-In AND~
219 274 1476 0 3 22
0 17 15 27
0
0 0 624 180
5 74F08
-18 -24 17 -16
3 U6D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
8186 0 0
2
43796 8
0
9 2-In AND~
219 273 1436 0 3 22
0 17 16 28
0
0 0 624 180
5 74F08
-18 -24 17 -16
3 U6C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
3754 0 0
2
43796 9
0
9 Inverter~
13 276 1395 0 2 22
0 17 29
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U8A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
8708 0 0
2
43796 10
0
9 2-In XOR~
219 271 1341 0 3 22
0 16 17 25
0
0 0 624 512
6 74LS86
-21 -24 21 -16
2 SD
2 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3338 0 0
2
43796 11
0
5 4071~
219 769 2522 0 3 22
0 58 62 20
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U17A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 15 0
1 U
5546 0 0
2
5.89917e-315 0
0
5 4071~
219 649 2567 0 3 22
0 64 63 62
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U18A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 16 0
1 U
3295 0 0
2
5.89917e-315 5.26354e-315
0
5 4071~
219 701 2480 0 3 22
0 59 65 58
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 17 0
1 U
4923 0 0
2
5.89917e-315 5.30499e-315
0
5 4081~
219 588 2400 0 3 22
0 18 34 66
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U25B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 20 0
1 U
3248 0 0
2
5.89917e-315 5.32571e-315
0
5 4071~
219 658 2377 0 3 22
0 67 66 19
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U20A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 34 0
1 U
3139 0 0
2
5.89917e-315 5.34643e-315
0
5 4081~
219 589 2348 0 3 22
0 18 35 67
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U25C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 20 0
1 U
3285 0 0
2
5.89917e-315 5.3568e-315
0
9 Inverter~
13 206 2289 0 2 22
0 18 41
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U21A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 35 0
1 U
336 0 0
2
5.89917e-315 5.36716e-315
0
9 Inverter~
13 253 2291 0 2 22
0 34 38
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U21B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 35 0
1 U
6582 0 0
2
5.89917e-315 5.37752e-315
0
9 Inverter~
13 300 2292 0 2 22
0 35 40
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U21C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 35 0
1 U
3546 0 0
2
5.89917e-315 5.38788e-315
0
9 Inverter~
13 346 2292 0 2 22
0 36 39
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U21D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 35 0
1 U
893 0 0
2
5.89917e-315 5.39306e-315
0
9 Inverter~
13 395 2291 0 2 22
0 24 61
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U21E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 35 0
1 U
8998 0 0
2
5.89917e-315 5.39824e-315
0
2 +V
167 163 2217 0 1 3
0 37
0
0 0 54256 0
2 5v
-8 -22 6 -14
2 V6
-8 -32 6 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5979 0 0
2
5.89917e-315 5.40342e-315
0
14 Logic Display~
6 797 2357 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.89917e-315 5.4086e-315
0
14 Logic Display~
6 857 2500 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
750 0 0
2
5.89917e-315 5.41378e-315
0
5 4073~
219 581 2499 0 4 22
0 41 34 35 65
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U37B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 32 0
1 U
849 0 0
2
5.89917e-315 5.41896e-315
0
5 4073~
219 582 2543 0 4 22
0 18 38 40 64
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U37C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 32 0
1 U
4693 0 0
2
5.89917e-315 5.42414e-315
0
5 4073~
219 582 2588 0 4 22
0 34 35 36 63
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U23A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 36 0
1 U
4775 0 0
2
5.89917e-315 5.42933e-315
0
5 4023~
219 581 2463 0 4 22
0 41 34 36 60
0
0 0 624 0
4 4023
-14 -28 14 -20
4 U38B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 33 0
1 U
9572 0 0
2
5.89917e-315 5.43192e-315
0
9 Inverter~
13 649 2472 0 2 22
0 60 59
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U21F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 35 0
1 U
3761 0 0
2
5.89917e-315 5.43451e-315
0
14 Logic Display~
6 834 2678 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6765 0 0
2
5.89917e-315 5.4371e-315
0
5 4071~
219 700 2698 0 3 22
0 55 54 21
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U20B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 34 0
1 U
7938 0 0
2
5.89917e-315 5.43969e-315
0
5 4071~
219 644 2664 0 3 22
0 57 56 55
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U20C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 34 0
1 U
55 0 0
2
5.89917e-315 5.44228e-315
0
5 4082~
219 573 2726 0 5 22
0 18 34 35 39 54
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U35B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 30 0
1 U
5610 0 0
2
5.89917e-315 5.44487e-315
0
5 4082~
219 572 2673 0 5 22
0 18 38 40 36 56
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U39A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 37 0
1 U
3322 0 0
2
5.89917e-315 5.44746e-315
0
5 4082~
219 574 2629 0 5 22
0 41 34 40 39 57
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U39B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 37 0
1 U
5914 0 0
2
5.89917e-315 5.45005e-315
0
14 Logic Display~
6 855 2801 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.89917e-315 5.45264e-315
0
5 4082~
219 571 2769 0 5 22
0 41 38 35 37 53
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U40A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 38 0
1 U
5830 0 0
2
5.89917e-315 5.45523e-315
0
5 4082~
219 571 2812 0 5 22
0 41 35 36 37 52
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U40B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 38 0
1 U
9153 0 0
2
5.89917e-315 5.45782e-315
0
5 4082~
219 570 2855 0 5 22
0 18 40 39 37 51
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U41A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 39 0
1 U
9220 0 0
2
5.89917e-315 5.46041e-315
0
5 4082~
219 569 2902 0 5 22
0 18 34 40 37 50
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U41B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 39 0
1 U
7901 0 0
2
5.89917e-315 5.463e-315
0
5 4071~
219 630 2786 0 3 22
0 53 52 48
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U20D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 34 0
1 U
4571 0 0
2
5.89917e-315 5.46559e-315
0
5 4071~
219 641 2870 0 3 22
0 51 50 49
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U42A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 40 0
1 U
7796 0 0
2
5.89917e-315 5.46818e-315
0
5 4071~
219 721 2821 0 3 22
0 48 49 22
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U42B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 40 0
1 U
3907 0 0
2
5.89917e-315 5.47077e-315
0
14 Logic Display~
6 855 2973 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4389 0 0
2
5.89917e-315 5.47207e-315
0
5 4071~
219 721 2994 0 3 22
0 42 43 23
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U42C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 40 0
1 U
7762 0 0
2
5.89917e-315 5.47336e-315
0
5 4071~
219 641 3043 0 3 22
0 45 44 43
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U42D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 40 0
1 U
6723 0 0
2
5.89917e-315 5.47466e-315
0
5 4071~
219 630 2959 0 3 22
0 47 46 42
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U43A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 41 0
1 U
6871 0 0
2
5.89917e-315 5.47595e-315
0
5 4082~
219 569 3075 0 5 22
0 38 35 36 37 44
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U44A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 42 0
1 U
4198 0 0
2
5.89917e-315 5.47725e-315
0
5 4082~
219 570 3028 0 5 22
0 18 38 40 39 45
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U44B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 42 0
1 U
970 0 0
2
5.89917e-315 5.47854e-315
0
5 4082~
219 571 2985 0 5 22
0 41 34 35 39 46
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U45A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 43 0
1 U
319 0 0
2
5.89917e-315 5.47984e-315
0
5 4082~
219 571 2942 0 5 22
0 41 38 36 37 47
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U45B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 43 0
1 U
3663 0 0
2
5.89917e-315 5.48113e-315
0
14 Logic Display~
6 848 3093 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3512 0 0
2
5.89917e-315 5.48243e-315
0
12 Hex Display~
7 1007 2287 0 18 19
10 20 19 144 145 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP8
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
7555 0 0
2
5.89917e-315 5.48372e-315
0
12 Hex Display~
7 1073 2286 0 18 19
10 24 23 22 21 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP9
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9776 0 0
2
5.89917e-315 5.48502e-315
0
5 4013~
219 880 1819 0 6 22
0 2 18 69 2 146 68
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U48B
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 46 0
1 U
6596 0 0
2
5.89917e-315 5.48631e-315
0
5 4013~
219 806 1818 0 6 22
0 2 34 69 2 147 76
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U48A
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 46 0
1 U
6750 0 0
2
5.89917e-315 5.48761e-315
0
5 4013~
219 730 1815 0 6 22
0 2 35 69 2 148 77
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U47B
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 45 0
1 U
9636 0 0
2
5.89917e-315 5.4889e-315
0
5 4013~
219 655 1819 0 6 22
0 2 36 69 2 149 78
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U47A
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 45 0
1 U
5369 0 0
2
5.89917e-315 5.4902e-315
0
7 Ground~
168 545 1674 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8555 0 0
2
5.89917e-315 5.49149e-315
0
7 Pulser~
4 490 1804 0 10 12
0 150 151 152 69 0 0 5 5 5
7
0
0 0 4656 0
0
2 V8
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4690 0 0
2
5.89917e-315 5.49279e-315
0
5 4013~
219 572 1820 0 6 22
0 2 24 69 2 153 71
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U46B
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 44 0
1 U
9145 0 0
2
5.89917e-315 5.49408e-315
0
9 2-In AND~
219 533 2047 0 3 22
0 71 79 70
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U6B
14 -20 35 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
5246 0 0
2
5.89917e-315 5.49538e-315
0
4 4008
219 565 1907 0 14 29
0 68 76 77 78 2 73 74 75 70
36 35 34 18 154
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U7
-8 -61 6 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9111 0 0
2
5.89917e-315 5.49667e-315
0
9 2-In AND~
219 226 2108 0 3 22
0 29 72 75
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U6A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6717 0 0
2
5.89917e-315 5.49797e-315
0
9 2-In AND~
219 282 2109 0 3 22
0 25 72 74
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 COUD
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3487 0 0
2
5.89917e-315 5.49926e-315
0
9 2-In AND~
219 347 2113 0 3 22
0 2 72 73
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 COUC
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
9604 0 0
2
5.89917e-315 5.50056e-315
0
9 2-In AND~
219 170 2105 0 3 22
0 26 72 79
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 COUB
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3921 0 0
2
5.89917e-315 5.50185e-315
0
9 2-In XOR~
219 479 2054 0 3 22
0 79 71 24
0
0 0 624 90
6 74LS86
-22 -24 20 -16
2 SC
-21 -25 -7 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 4 0
1 U
8146 0 0
2
5.89917e-315 5.50315e-315
0
7 Ground~
168 302 1902 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4506 0 0
2
5.89917e-315 5.50444e-315
0
2 +V
167 402 187 0 1 3
0 87
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5386 0 0
2
5.89917e-315 5.50574e-315
0
9 CA 7-Seg~
184 403 233 0 18 19
10 86 85 84 83 82 81 80 155 87
0 0 2 0 0 2 0 2 1
0
0 0 21088 0
8 YELLOWCA
6 -41 62 -33
4 DADO
33 -4 61 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7847 0 0
2
5.89917e-315 5.50703e-315
0
12 Hex Display~
7 471 108 0 18 19
10 20 19 156 157 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP5
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9261 0 0
2
43796 12
0
12 Hex Display~
7 504 108 0 18 19
10 24 23 22 21 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8231 0 0
2
43796 13
0
12 Hex Display~
7 321 113 0 18 19
10 13 12 11 10 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP6
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3756 0 0
2
43796 14
0
12 Hex Display~
7 288 113 0 18 19
10 9 8 158 159 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
6760 0 0
2
43796 15
0
2 +V
167 97 569 0 1 3
0 89
0
0 0 54256 0
2 5V
-8 -20 6 -12
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
351 0 0
2
43796 16
0
7 Ground~
168 611 680 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
5352 0 0
2
5.89917e-315 5.50833e-315
0
5 4013~
219 1420 575 0 6 22
0 2 30 94 2 160 90
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U14B
17 -61 45 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 8 0
1 U
485 0 0
2
5.89917e-315 5.50963e-315
0
14 NO PushButton~
191 72 184 0 2 5
0 89 72
0
0 0 4720 0
0
5 Jogar
-13 -26 22 -18
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
452 0 0
2
5.89917e-315 5.51092e-315
0
9 2-In AND~
219 843 825 0 3 22
0 98 17 99
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 COUT
11 -20 39 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
643 0 0
2
5.89917e-315 5.51222e-315
0
9 2-In XOR~
219 788 832 0 3 22
0 17 98 13
0
0 0 624 90
6 74LS86
-22 -24 20 -16
2 S0
-21 -25 -7 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 102
65 0 0 0 4 1 4 0
1 U
5563 0 0
2
5.89917e-315 5.51286e-315
0
12 Hex Display~
7 644 478 0 18 19
10 98 97 96 95 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
934 0 0
2
5.89917e-315 5.51351e-315
0
5 4071~
219 1587 1272 0 3 22
0 119 122 9
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U30B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 25 0
1 U
3240 0 0
2
5.89917e-315 5.51416e-315
0
5 4071~
219 1467 1317 0 3 22
0 124 123 122
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U30A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 25 0
1 U
3233 0 0
2
5.89917e-315 5.51481e-315
0
5 4071~
219 1519 1230 0 3 22
0 120 125 119
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U24D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 19 0
1 U
3635 0 0
2
5.89917e-315 5.51545e-315
0
5 4081~
219 1406 1150 0 3 22
0 30 91 126
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U25A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 20 0
1 U
3547 0 0
2
5.89917e-315 5.5161e-315
0
5 4071~
219 1476 1127 0 3 22
0 127 126 8
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U24A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 19 0
1 U
483 0 0
2
5.89917e-315 5.51675e-315
0
5 4081~
219 1407 1098 0 3 22
0 30 92 127
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 18 0
1 U
6126 0 0
2
5.89917e-315 5.5174e-315
0
9 Inverter~
13 1024 1039 0 2 22
0 30 31
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U36A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 31 0
1 U
7368 0 0
2
5.89917e-315 5.51804e-315
0
9 Inverter~
13 1071 1041 0 2 22
0 91 100
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U36B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 31 0
1 U
3925 0 0
2
5.89917e-315 5.51869e-315
0
9 Inverter~
13 1118 1042 0 2 22
0 92 102
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U36C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 31 0
1 U
6187 0 0
2
5.89917e-315 5.51934e-315
0
9 Inverter~
13 1164 1042 0 2 22
0 93 101
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U36D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 31 0
1 U
5866 0 0
2
5.89917e-315 5.51999e-315
0
9 Inverter~
13 1213 1041 0 2 22
0 13 32
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U36E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 31 0
1 U
6650 0 0
2
5.89917e-315 5.52063e-315
0
2 +V
167 981 967 0 1 3
0 33
0
0 0 54256 0
2 5v
-8 -22 6 -14
3 V16
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8814 0 0
2
5.89917e-315 5.52128e-315
0
14 Logic Display~
6 1615 1107 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4714 0 0
2
5.89917e-315 5.52193e-315
0
14 Logic Display~
6 1675 1250 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9875 0 0
2
5.89917e-315 5.52258e-315
0
5 4073~
219 1399 1249 0 4 22
0 31 91 92 125
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U28B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 23 0
1 U
8220 0 0
2
5.89917e-315 5.52322e-315
0
5 4073~
219 1400 1293 0 4 22
0 30 100 102 124
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U28C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 23 0
1 U
3691 0 0
2
5.89917e-315 5.52387e-315
0
5 4073~
219 1400 1338 0 4 22
0 91 92 93 123
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U37A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 32 0
1 U
5196 0 0
2
5.89917e-315 5.52452e-315
0
5 4023~
219 1399 1213 0 4 22
0 31 91 93 121
0
0 0 624 0
4 4023
-14 -28 14 -20
4 U38A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 33 0
1 U
6182 0 0
2
5.89917e-315 5.52517e-315
0
9 Inverter~
13 1467 1222 0 2 22
0 121 120
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U36F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 31 0
1 U
6326 0 0
2
5.89917e-315 5.52581e-315
0
14 Logic Display~
6 1652 1428 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3247 0 0
2
5.89917e-315 5.52646e-315
0
5 4071~
219 1518 1448 0 3 22
0 116 115 10
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U24C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 19 0
1 U
5235 0 0
2
5.89917e-315 5.52711e-315
0
5 4071~
219 1462 1414 0 3 22
0 118 117 116
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U24B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 19 0
1 U
9260 0 0
2
5.89917e-315 5.52776e-315
0
5 4082~
219 1391 1476 0 5 22
0 30 91 92 101 115
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U27A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 22 0
1 U
583 0 0
2
5.89917e-315 5.52841e-315
0
5 4082~
219 1390 1423 0 5 22
0 30 100 102 93 117
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U26B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 21 0
1 U
3471 0 0
2
5.89917e-315 5.52905e-315
0
5 4082~
219 1392 1379 0 5 22
0 31 91 102 101 118
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U26A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 21 0
1 U
7124 0 0
2
5.89917e-315 5.5297e-315
0
14 Logic Display~
6 1673 1551 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6160 0 0
2
5.89917e-315 5.53035e-315
0
5 4082~
219 1389 1519 0 5 22
0 31 100 92 33 114
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U29B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 24 0
1 U
4732 0 0
2
5.89917e-315 5.531e-315
0
5 4082~
219 1389 1562 0 5 22
0 31 92 93 33 113
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U31A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 26 0
1 U
8836 0 0
2
5.89917e-315 5.53164e-315
0
5 4082~
219 1388 1605 0 5 22
0 30 102 101 33 112
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U31B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 26 0
1 U
3346 0 0
2
5.89917e-315 5.53229e-315
0
5 4082~
219 1387 1652 0 5 22
0 30 91 102 33 111
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U32A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 27 0
1 U
8546 0 0
2
5.89917e-315 5.53294e-315
0
5 4071~
219 1448 1536 0 3 22
0 114 113 109
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U30C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 25 0
1 U
8607 0 0
2
5.89917e-315 5.53359e-315
0
5 4071~
219 1459 1620 0 3 22
0 112 111 110
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U30D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 25 0
1 U
5781 0 0
2
5.89917e-315 5.53423e-315
0
5 4071~
219 1539 1571 0 3 22
0 109 110 11
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U33A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 28 0
1 U
6991 0 0
2
5.89917e-315 5.53488e-315
0
14 Logic Display~
6 1673 1723 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9631 0 0
2
5.89917e-315 5.53553e-315
0
5 4071~
219 1539 1744 0 3 22
0 103 104 12
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U33B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 28 0
1 U
8381 0 0
2
5.89917e-315 5.53618e-315
0
5 4071~
219 1459 1793 0 3 22
0 106 105 104
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U33C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 28 0
1 U
6697 0 0
2
5.89917e-315 5.53682e-315
0
5 4071~
219 1448 1709 0 3 22
0 108 107 103
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U33D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 28 0
1 U
3463 0 0
2
5.89917e-315 5.53747e-315
0
5 4082~
219 1387 1825 0 5 22
0 100 92 93 30 105
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U32B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 27 0
1 U
9605 0 0
2
5.89917e-315 5.53812e-315
0
5 4082~
219 1388 1778 0 5 22
0 30 100 102 101 106
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U34A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 29 0
1 U
936 0 0
2
5.89917e-315 5.53877e-315
0
5 4082~
219 1389 1735 0 5 22
0 31 91 92 101 107
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U34B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 29 0
1 U
9813 0 0
2
5.89917e-315 5.53941e-315
0
5 4082~
219 1389 1692 0 5 22
0 31 100 93 33 108
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U35A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 30 0
1 U
5286 0 0
2
5.89917e-315 5.54006e-315
0
14 Logic Display~
6 1666 1843 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9179 0 0
2
5.89917e-315 5.54071e-315
0
7 Ground~
168 826 415 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3718 0 0
2
43796 17
0
5 4013~
219 1290 571 0 6 22
0 2 91 94 2 161 95
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U14A
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 8 0
1 U
4375 0 0
2
43796 18
0
5 4013~
219 1143 575 0 6 22
0 2 92 94 2 162 96
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U12B
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 7 0
1 U
3616 0 0
2
43796 19
0
5 4013~
219 1005 575 0 6 22
0 2 93 94 2 163 97
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U12A
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 7 0
1 U
7808 0 0
2
43796 20
0
14 Logic Display~
6 820 586 0 1 2
10 94
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7498 0 0
2
43796 21
0
5 4013~
219 862 563 0 6 22
0 2 13 94 2 164 98
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U9B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
9736 0 0
2
43796 22
0
4 4008
219 876 685 0 14 29
0 90 95 96 97 2 2 15 16 99
93 92 91 30 165
0
0 0 4848 0
4 4008
-14 -60 14 -52
3 U10
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9454 0 0
2
43796 23
0
7 Pulser~
4 763 557 0 10 12
0 166 167 168 94 0 0 5 5 5
7
0
0 0 4656 0
0
2 V7
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4639 0 0
2
43796 24
0
9 2-In AND~
219 479 883 0 3 22
0 133 72 17
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U5D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3831 0 0
2
43796 25
0
9 2-In AND~
219 656 891 0 3 22
0 130 72 2
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U5C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3538 0 0
2
43796 26
0
9 2-In AND~
219 591 887 0 3 22
0 131 72 15
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U5B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5949 0 0
2
43796 27
0
9 2-In AND~
219 535 886 0 3 22
0 132 72 16
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U5A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7130 0 0
2
43796 28
0
10 2-In XNOR~
219 409 1221 0 3 22
0 2 133 134
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4D
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
4115 0 0
2
43796 29
0
10 2-In XNOR~
219 410 1184 0 3 22
0 128 132 135
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4C
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3197 0 0
2
43796 30
0
10 2-In XNOR~
219 411 1143 0 3 22
0 128 131 136
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4B
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
813 0 0
2
43796 31
0
10 2-In XNOR~
219 411 1106 0 3 22
0 2 130 137
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4A
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3396 0 0
2
43796 32
0
5 7422~
219 329 1153 0 5 22
0 134 136 135 137 138
0
0 0 624 180
6 74LS22
-21 -28 21 -20
3 U3A
-8 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
6348 0 0
2
43796 33
0
7 Ground~
168 329 1044 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
583 0 0
2
43796 34
0
14 Logic Display~
6 135 900 0 1 2
10 139
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
922 0 0
2
43796 35
0
7 Pulser~
4 60 971 0 10 12
0 169 170 139 171 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4442 0 0
2
43796 36
0
6 74LS47
187 663 1026 0 14 29
0 130 131 132 133 172 173 80 81 82
83 84 85 86 174
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5893 0 0
2
43796 37
0
7 74LS190
134 380 980 0 14 29
0 72 139 138 129 2 2 2 128 175
176 130 131 132 133
0
0 0 4848 0
6 74F190
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3814 0 0
2
43796 38
0
7 Ground~
168 640 1135 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3637 0 0
2
43796 39
0
2 +V
167 596 1165 0 1 3
0 128
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6890 0 0
2
43796 40
0
7 Ground~
168 339 723 0 1 3
0 2
0
0 0 53360 180
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3933 0 0
2
43796 41
0
9 Resistor~
219 215 754 0 4 5
0 72 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3432 0 0
2
43796 42
0
418
1 14 3 0 0 8320 0 2 7 0 0 5
496 217
496 254
1636 254
1636 724
1542 724
0 0 2 0 0 4096 0 0 0 370 373 2
944 581
944 411
1 0 4 0 0 0 0 3 0 0 4 2
275 225
275 225
13 0 4 0 0 12416 0 7 0 0 0 5
1542 715
1596 715
1596 325
275 325
275 221
9 12 5 0 0 8320 0 7 6 0 0 4
1542 661
1575 661
1575 812
1542 812
10 13 6 0 0 8320 0 7 6 0 0 4
1542 670
1564 670
1564 821
1542 821
11 14 7 0 0 8320 0 7 6 0 0 4
1542 679
1556 679
1556 830
1542 830
3 0 8 0 0 8192 0 7 0 0 266 3
1478 679
1341 679
1341 13
4 0 9 0 0 8192 0 7 0 0 267 3
1478 688
1356 688
1356 9
0 1 10 0 0 4096 0 0 6 275 0 3
1400 51
1400 767
1478 767
2 0 11 0 0 8192 0 6 0 0 276 3
1478 776
1391 776
1391 46
3 0 12 0 0 8192 0 6 0 0 277 3
1478 785
1380 785
1380 44
0 4 13 0 0 4096 0 0 6 278 0 3
1365 40
1365 794
1478 794
0 4 2 0 0 0 0 0 82 368 0 2
1290 581
1420 581
8 0 14 0 0 4096 0 6 0 0 22 2
1478 830
1350 830
7 0 2 0 0 0 0 6 0 0 24 2
1478 821
1374 821
6 0 2 0 0 0 0 6 0 0 24 2
1478 812
1374 812
5 0 2 0 0 0 0 6 0 0 24 2
1478 803
1374 803
8 0 2 0 0 0 0 7 0 0 24 2
1478 724
1374 724
7 0 14 0 0 0 0 7 0 0 22 2
1478 715
1350 715
0 0 2 0 0 0 0 0 0 24 23 2
1374 705
1470 705
0 1 14 0 0 4224 0 0 4 0 0 2
1350 665
1350 837
5 6 2 0 0 0 0 7 7 0 0 4
1478 697
1470 697
1470 706
1478 706
2 1 2 0 0 16384 0 7 5 0 0 5
1478 670
1470 670
1470 666
1374 666
1374 846
1 0 2 0 0 0 0 7 0 0 24 3
1478 661
1470 661
1470 666
0 0 2 0 0 0 0 0 0 25 25 4
1470 665
1469 665
1469 665
1470 665
0 0 2 0 0 0 0 0 0 201 35 2
108 1337
108 1323
2 0 15 0 0 8320 0 11 0 0 244 5
292 1467
785 1467
785 894
695 894
695 703
2 0 16 0 0 4096 0 12 0 0 34 3
291 1427
745 1427
745 1332
1 0 17 0 0 4096 0 11 0 0 31 3
292 1485
757 1485
757 1445
1 0 17 0 0 4096 0 12 0 0 32 3
291 1445
757 1445
757 1395
1 0 17 0 0 0 0 13 0 0 33 3
297 1395
757 1395
757 1350
2 0 17 0 0 8320 0 14 0 0 256 3
293 1350
757 1350
757 859
1 0 16 0 0 8320 0 14 0 0 245 3
293 1332
745 1332
745 712
4 1 2 0 0 0 0 9 8 0 0 4
66 1323
133 1323
133 1295
160 1295
0 0 2 0 0 0 0 0 0 243 37 2
780 694
780 685
5 1 2 0 0 12416 0 135 8 0 0 4
844 685
773 685
773 1295
160 1295
1 0 18 0 0 4096 0 43 0 0 72 2
546 2842
237 2842
0 2 19 0 0 8320 0 0 76 69 0 5
1010 2370
1861 2370
1861 164
474 164
474 132
1 0 20 0 0 12416 0 76 0 0 70 5
480 132
480 159
1851 159
1851 2363
1016 2363
4 0 21 0 0 12416 0 77 0 0 65 5
495 132
495 152
1814 152
1814 2346
1064 2346
0 3 22 0 0 8320 0 0 77 43 0 4
1820 1215
1820 146
501 146
501 132
0 0 22 0 0 0 0 0 0 66 42 3
1070 2335
1820 2335
1820 1209
2 0 23 0 0 12416 0 77 0 0 67 5
507 132
507 140
1825 140
1825 2327
1076 2327
1 0 24 0 0 8320 0 77 0 0 68 4
513 132
1835 132
1835 2319
1082 2319
3 3 25 0 0 4096 0 14 9 0 0 3
244 1341
72 1341
72 1323
3 1 26 0 0 8192 0 10 9 0 0 3
175 1455
84 1455
84 1323
2 3 27 0 0 4224 0 10 11 0 0 4
221 1464
241 1464
241 1476
247 1476
1 3 28 0 0 4224 0 10 12 0 0 4
221 1446
240 1446
240 1436
246 1436
2 2 29 0 0 8192 0 9 13 0 0 3
78 1323
78 1395
261 1395
1 0 30 0 0 4096 0 115 0 0 240 2
1364 1592
1053 1592
0 0 24 0 0 0 0 0 0 53 83 3
482 2015
418 2015
418 2275
2 3 24 0 0 0 0 65 72 0 0 7
548 1784
529 1784
529 1758
446 1758
446 1987
482 1987
482 2024
0 0 31 0 0 4096 0 0 0 289 0 2
1027 1722
1027 1990
4 0 2 0 0 0 0 59 0 0 195 2
880 1825
880 1857
4 0 2 0 0 0 0 60 0 0 195 2
806 1824
806 1857
4 0 2 0 0 0 0 62 0 0 195 2
655 1825
655 1857
4 0 2 0 0 0 0 61 0 0 195 2
730 1821
730 1857
2 0 32 0 0 4224 0 97 0 0 0 2
1216 1059
1216 1966
0 0 33 0 0 4096 0 0 0 290 0 2
983 1706
983 1980
0 0 18 0 0 8320 0 0 0 180 77 6
799 1889
799 2174
234 2174
234 2227
235 2227
235 2272
0 0 34 0 0 8320 0 0 0 181 157 4
768 1897
768 2190
278 2190
278 2275
0 0 35 0 0 8320 0 0 0 182 158 4
698 1907
698 2217
325 2217
325 2276
0 0 36 0 0 4224 0 0 0 183 155 4
610 1916
610 2232
368 2232
368 2274
4 1 21 0 0 0 0 58 34 0 0 3
1064 2310
1064 2696
834 2696
1 3 22 0 0 0 0 40 58 0 0 3
855 2819
1070 2819
1070 2310
2 0 23 0 0 0 0 58 0 0 100 3
1076 2310
1076 2993
855 2993
1 1 24 0 0 0 0 56 58 0 0 3
848 3111
1082 3111
1082 2310
1 2 19 0 0 0 0 27 57 0 0 3
797 2375
1010 2375
1010 2311
1 1 20 0 0 0 0 28 57 0 0 3
857 2518
1016 2518
1016 2311
1 0 18 0 0 0 0 53 0 0 72 3
546 3015
237 3015
237 2889
1 0 18 0 0 0 0 44 0 0 73 3
545 2889
237 2889
237 2713
1 0 18 0 0 0 0 37 0 0 74 3
549 2713
237 2713
237 2660
1 0 18 0 0 0 0 38 0 0 75 3
548 2660
237 2660
237 2534
1 0 18 0 0 0 0 30 0 0 76 3
558 2534
235 2534
235 2391
1 0 18 0 0 0 0 18 0 0 77 3
564 2391
235 2391
235 2339
1 1 18 0 0 0 0 20 21 0 0 4
565 2339
235 2339
235 2271
209 2271
0 0 36 0 0 0 0 0 0 85 0 2
372 3080
372 3248
0 0 35 0 0 0 0 0 0 86 0 2
325 3071
325 3250
0 0 34 0 0 0 0 0 0 81 0 2
281 2981
281 3247
0 0 34 0 0 0 0 0 0 82 93 2
281 2898
281 2981
0 0 34 0 0 0 0 0 0 132 111 2
281 2722
281 2898
1 1 24 0 0 0 0 56 25 0 0 4
848 3111
418 3111
418 2273
398 2273
4 0 37 0 0 4096 0 52 0 0 165 2
545 3089
163 3089
3 0 36 0 0 0 0 52 0 0 96 3
545 3080
369 3080
369 2947
2 0 35 0 0 0 0 52 0 0 92 3
545 3071
325 3071
325 2990
1 0 38 0 0 4096 0 52 0 0 170 2
545 3062
256 3062
4 0 39 0 0 4096 0 53 0 0 168 2
546 3042
349 3042
3 0 40 0 0 4096 0 53 0 0 169 2
546 3033
303 3033
2 0 38 0 0 4096 0 53 0 0 170 2
546 3024
256 3024
4 0 39 0 0 4096 0 54 0 0 168 2
547 2999
349 2999
3 0 35 0 0 0 0 54 0 0 117 3
547 2990
325 2990
325 2808
2 0 34 0 0 0 0 54 0 0 0 2
547 2981
278 2981
1 0 41 0 0 4096 0 54 0 0 171 2
547 2972
209 2972
4 0 37 0 0 4096 0 55 0 0 165 2
547 2956
163 2956
3 0 36 0 0 0 0 55 0 0 116 3
547 2947
369 2947
369 2817
2 0 38 0 0 4096 0 55 0 0 170 2
547 2938
256 2938
1 0 41 0 0 0 0 55 0 0 171 2
547 2929
209 2929
3 0 23 0 0 0 0 49 0 0 100 2
754 2994
754 2993
1 3 23 0 0 0 0 48 0 0 0 3
855 2991
855 2993
749 2993
0 3 36 0 0 0 0 0 52 0 0 3
553 3081
553 3080
545 3080
3 1 42 0 0 4224 0 51 49 0 0 4
663 2959
700 2959
700 2985
708 2985
3 2 43 0 0 8320 0 50 49 0 0 4
674 3043
700 3043
700 3003
708 3003
5 2 44 0 0 4224 0 52 50 0 0 4
590 3075
620 3075
620 3052
628 3052
5 1 45 0 0 4224 0 53 50 0 0 4
591 3028
620 3028
620 3034
628 3034
5 2 46 0 0 4224 0 54 51 0 0 4
592 2985
609 2985
609 2968
617 2968
5 1 47 0 0 4224 0 55 51 0 0 4
592 2942
609 2942
609 2950
617 2950
3 0 35 0 0 0 0 41 0 0 131 3
547 2774
325 2774
325 2731
4 0 37 0 0 0 0 44 0 0 165 2
545 2916
163 2916
3 0 40 0 0 0 0 44 0 0 169 2
545 2907
303 2907
2 0 34 0 0 0 0 44 0 0 0 2
545 2898
278 2898
4 0 37 0 0 0 0 43 0 0 165 2
546 2869
163 2869
3 0 39 0 0 0 0 43 0 0 168 2
546 2860
349 2860
2 0 40 0 0 0 0 43 0 0 169 2
546 2851
303 2851
4 0 37 0 0 0 0 42 0 0 165 2
547 2826
163 2826
3 0 36 0 0 0 0 42 0 0 133 3
547 2817
368 2817
368 2687
2 0 35 0 0 0 0 42 0 0 108 3
547 2808
325 2808
325 2774
1 0 41 0 0 0 0 42 0 0 171 2
547 2799
209 2799
4 0 37 0 0 0 0 41 0 0 165 2
547 2783
163 2783
2 0 38 0 0 0 0 41 0 0 170 2
547 2765
256 2765
1 0 41 0 0 0 0 41 0 0 171 2
547 2756
209 2756
3 0 22 0 0 0 0 47 0 0 123 2
754 2821
754 2821
1 3 22 0 0 0 0 40 0 0 0 3
855 2819
855 2821
749 2821
3 1 48 0 0 4224 0 45 47 0 0 4
663 2786
700 2786
700 2812
708 2812
3 2 49 0 0 8320 0 46 47 0 0 4
674 2870
700 2870
700 2830
708 2830
5 2 50 0 0 4224 0 44 46 0 0 4
590 2902
620 2902
620 2879
628 2879
5 1 51 0 0 4224 0 43 46 0 0 4
591 2855
620 2855
620 2861
628 2861
5 2 52 0 0 4224 0 42 45 0 0 4
592 2812
609 2812
609 2795
617 2795
5 1 53 0 0 4224 0 41 45 0 0 4
592 2769
609 2769
609 2777
617 2777
4 0 39 0 0 4096 0 37 0 0 168 2
549 2740
349 2740
3 0 35 0 0 0 0 37 0 0 149 3
549 2731
325 2731
325 2588
2 0 34 0 0 0 0 37 0 0 138 3
549 2722
279 2722
279 2625
4 0 36 0 0 0 0 38 0 0 148 3
548 2687
368 2687
368 2597
3 0 40 0 0 4096 0 38 0 0 169 2
548 2678
303 2678
2 0 38 0 0 4096 0 38 0 0 170 2
548 2669
256 2669
4 0 39 0 0 4096 0 39 0 0 168 2
550 2643
349 2643
3 0 40 0 0 4096 0 39 0 0 169 2
550 2634
303 2634
2 0 34 0 0 0 0 39 0 0 150 3
550 2625
279 2625
279 2579
1 0 41 0 0 4096 0 39 0 0 171 2
550 2616
209 2616
3 0 21 0 0 0 0 35 0 0 141 2
733 2698
733 2698
1 3 21 0 0 0 0 34 0 0 0 3
834 2696
834 2698
728 2698
5 2 54 0 0 4224 0 37 35 0 0 4
594 2726
679 2726
679 2707
687 2707
1 3 55 0 0 8320 0 35 36 0 0 3
687 2689
677 2689
677 2664
5 2 56 0 0 4224 0 38 36 0 0 2
593 2673
631 2673
5 1 57 0 0 4224 0 39 36 0 0 4
595 2629
623 2629
623 2655
631 2655
1 0 41 0 0 4096 0 29 0 0 171 2
557 2490
209 2490
1 0 41 0 0 0 0 32 0 0 171 2
557 2454
209 2454
3 0 36 0 0 0 0 31 0 0 155 3
558 2597
368 2597
368 2472
2 0 35 0 0 0 0 31 0 0 153 3
558 2588
325 2588
325 2508
1 0 34 0 0 0 0 31 0 0 154 3
558 2579
279 2579
279 2499
3 0 40 0 0 4096 0 30 0 0 169 2
558 2552
303 2552
2 0 38 0 0 4096 0 30 0 0 170 2
558 2543
256 2543
3 0 35 0 0 0 0 29 0 0 158 3
557 2508
325 2508
325 2357
2 0 34 0 0 0 0 29 0 0 156 3
557 2499
278 2499
278 2463
3 1 36 0 0 0 0 32 24 0 0 4
557 2472
368 2472
368 2274
349 2274
2 0 34 0 0 0 0 32 0 0 157 3
557 2463
278 2463
278 2409
2 1 34 0 0 0 0 18 22 0 0 4
564 2409
278 2409
278 2273
256 2273
2 1 35 0 0 0 0 20 23 0 0 4
565 2357
325 2357
325 2274
303 2274
3 1 20 0 0 0 0 15 28 0 0 3
802 2522
857 2522
857 2518
3 1 58 0 0 4224 0 17 15 0 0 3
734 2480
734 2513
756 2513
2 1 59 0 0 8320 0 33 17 0 0 3
670 2472
670 2471
688 2471
4 0 60 0 0 0 0 32 0 0 176 2
608 2463
608 2463
2 0 39 0 0 0 0 24 0 0 168 2
349 2310
349 2310
1 3 19 0 0 0 0 27 19 0 0 3
797 2375
797 2377
691 2377
1 0 37 0 0 4224 0 26 0 0 0 2
163 2226
163 3251
2 0 61 0 0 4224 0 25 0 0 0 2
398 2309
398 3257
0 2 61 0 0 0 0 0 25 0 0 3
401 2308
401 2309
398 2309
0 0 39 0 0 4224 0 0 0 0 0 2
349 2301
349 3250
2 0 40 0 0 4224 0 23 0 0 0 2
303 2310
303 3256
2 0 38 0 0 4224 0 22 0 0 0 2
256 2309
256 3249
2 0 41 0 0 4224 0 21 0 0 0 2
209 2307
209 3251
3 2 62 0 0 12416 0 16 15 0 0 4
682 2567
703 2567
703 2531
756 2531
4 2 63 0 0 12416 0 31 16 0 0 6
603 2588
601 2588
601 2588
628 2588
628 2576
636 2576
4 1 64 0 0 4224 0 30 16 0 0 4
603 2543
628 2543
628 2558
636 2558
4 2 65 0 0 12416 0 29 17 0 0 4
602 2499
626 2499
626 2489
688 2489
0 1 60 0 0 4224 0 0 33 0 0 5
602 2463
626 2463
626 2471
634 2471
634 2472
2 3 66 0 0 4224 0 19 18 0 0 4
645 2386
608 2386
608 2400
609 2400
1 3 67 0 0 4224 0 19 20 0 0 3
645 2368
610 2368
610 2348
6 1 68 0 0 12416 0 59 67 0 0 6
904 1783
915 1783
915 1701
365 1701
365 1871
533 1871
13 2 18 0 0 0 0 67 59 0 0 4
597 1889
848 1889
848 1783
856 1783
2 12 34 0 0 0 0 60 67 0 0 4
782 1782
768 1782
768 1898
597 1898
11 2 35 0 0 0 0 67 61 0 0 4
597 1907
698 1907
698 1779
706 1779
2 10 36 0 0 0 0 62 67 0 0 3
631 1783
631 1916
597 1916
1 0 2 0 0 0 0 59 0 0 195 2
880 1762
880 1696
1 0 2 0 0 0 0 60 0 0 197 2
806 1761
806 1696
1 0 2 0 0 0 0 61 0 0 197 2
730 1758
730 1696
1 0 2 0 0 0 0 62 0 0 197 4
655 1762
655 1717
656 1717
656 1696
3 0 69 0 0 4096 0 59 0 0 198 2
856 1801
856 1838
3 0 69 0 0 4096 0 60 0 0 198 2
782 1800
782 1838
3 0 69 0 0 4096 0 61 0 0 198 2
706 1797
706 1838
3 0 69 0 0 0 0 62 0 0 198 3
631 1801
617 1801
617 1838
4 0 69 0 0 0 0 64 0 0 198 3
520 1804
520 1802
538 1802
4 0 30 0 0 0 0 124 0 0 240 2
1363 1839
1053 1839
0 0 2 0 0 0 0 0 0 195 195 4
970 1806
974 1806
974 1807
970 1807
4 0 2 0 0 0 0 65 0 0 197 5
572 1826
572 1857
970 1857
970 1696
857 1696
1 0 2 0 0 0 0 65 0 0 197 2
572 1763
572 1696
1 0 2 0 0 0 0 63 0 0 195 4
545 1668
572 1668
572 1696
861 1696
3 0 69 0 0 12416 0 65 0 0 0 4
548 1802
538 1802
538 1838
931 1838
9 3 70 0 0 8320 0 67 66 0 0 3
533 1943
532 1943
532 2023
2 1 71 0 0 20480 0 72 66 0 0 7
491 2073
492 2073
492 2072
491 2072
491 2090
523 2090
523 2068
1 0 2 0 0 0 0 70 0 0 0 5
337 2134
321 2134
321 1686
108 1686
108 1332
1 0 25 0 0 8320 0 69 0 0 46 5
272 2130
258 2130
258 1662
118 1662
118 1341
1 0 29 0 0 8320 0 68 0 0 50 5
216 2129
200 2129
200 1639
128 1639
128 1395
1 0 26 0 0 8320 0 71 0 0 47 3
160 2126
147 2126
147 1455
0 0 72 0 0 4224 0 0 0 232 216 2
27 754
27 2141
5 1 2 0 0 0 0 67 73 0 0 5
533 1907
337 1907
337 1889
302 1889
302 1896
3 6 73 0 0 8320 0 70 67 0 0 3
346 2089
346 1916
533 1916
3 7 74 0 0 8320 0 69 67 0 0 3
281 2085
281 1925
533 1925
3 8 75 0 0 8320 0 68 67 0 0 3
225 2084
225 1934
533 1934
6 2 76 0 0 8320 0 60 67 0 0 5
830 1782
830 1709
371 1709
371 1880
533 1880
6 3 77 0 0 8320 0 61 67 0 0 5
754 1779
754 1719
382 1719
382 1889
533 1889
6 4 78 0 0 8320 0 62 67 0 0 5
679 1783
679 1737
392 1737
392 1898
533 1898
6 0 71 0 0 16512 0 65 0 0 200 7
596 1784
601 1784
601 1728
404 1728
404 2072
491 2072
491 2073
3 0 79 0 0 4224 0 71 0 0 215 2
169 2081
473 2081
1 2 79 0 0 0 0 72 66 0 0 4
473 2073
473 2096
541 2096
541 2068
0 0 72 0 0 0 0 0 0 219 0 2
179 2141
21 2141
2 2 72 0 0 0 0 69 70 0 0 4
290 2130
290 2141
355 2141
355 2134
2 0 72 0 0 0 0 68 0 0 217 3
234 2129
234 2141
290 2141
2 0 72 0 0 0 0 71 0 0 218 3
178 2126
178 2141
234 2141
7 7 80 0 0 4224 0 75 149 0 0 5
418 269
418 919
739 919
739 990
701 990
6 8 81 0 0 4224 0 75 149 0 0 5
412 269
412 919
734 919
734 999
701 999
5 9 82 0 0 4224 0 75 149 0 0 5
406 269
406 919
729 919
729 1008
701 1008
4 10 83 0 0 4224 0 75 149 0 0 5
400 269
400 919
724 919
724 1017
701 1017
3 11 84 0 0 4224 0 75 149 0 0 5
394 269
394 919
719 919
719 1026
701 1026
2 12 85 0 0 4224 0 75 149 0 0 5
388 269
388 924
714 924
714 1035
701 1035
1 13 86 0 0 4224 0 75 149 0 0 5
382 269
382 929
709 929
709 1044
701 1044
1 0 87 0 0 4096 0 74 0 0 229 2
402 196
402 197
0 0 88 0 0 4224 0 0 0 0 0 3
140 1419
140 1417
139 1417
9 0 87 0 0 8320 0 75 0 0 0 5
403 197
402 197
402 195
403 195
403 194
1 1 89 0 0 16512 0 83 80 0 0 6
89 192
103 192
103 144
27 144
27 578
97 578
1 0 72 0 0 0 0 154 0 0 386 4
197 754
197 919
337 919
337 917
2 1 72 0 0 0 0 83 154 0 0 4
55 192
19 192
19 754
197 754
1 0 30 0 0 0 0 125 0 0 240 2
1364 1765
1053 1765
1 0 30 0 0 0 0 116 0 0 240 2
1363 1639
1053 1639
1 0 30 0 0 4096 0 109 0 0 240 2
1367 1463
1053 1463
1 0 30 0 0 0 0 110 0 0 240 2
1366 1410
1053 1410
1 0 30 0 0 4096 0 102 0 0 240 2
1376 1284
1053 1284
1 0 30 0 0 4096 0 90 0 0 240 2
1382 1141
1053 1141
1 0 30 0 0 4096 0 92 0 0 240 2
1383 1089
1053 1089
0 0 30 0 0 4224 0 0 0 257 0 2
1053 1020
1053 1998
1 0 2 0 0 0 0 82 0 0 371 3
1420 518
1420 411
1290 411
6 1 90 0 0 12416 0 82 135 0 0 6
1444 539
1449 539
1449 449
668 449
668 649
844 649
3 6 2 0 0 0 0 138 135 0 0 3
655 867
655 694
844 694
3 7 15 0 0 0 0 139 135 0 0 3
590 863
590 703
844 703
3 8 16 0 0 0 0 140 135 0 0 3
534 862
534 712
844 712
2 0 13 0 0 0 0 134 0 0 261 5
838 527
729 527
729 781
756 781
756 798
0 13 30 0 0 0 0 0 135 257 0 2
974 667
908 667
0 12 91 0 0 4096 0 0 135 258 0 2
947 676
908 676
0 11 92 0 0 4096 0 0 135 259 0 2
934 685
908 685
0 10 93 0 0 4096 0 0 135 260 0 2
919 694
908 694
0 3 94 0 0 4096 0 0 82 377 0 4
1209 616
1364 616
1364 557
1396 557
0 2 95 0 0 8192 0 0 135 268 0 3
680 551
680 658
844 658
0 3 96 0 0 8192 0 0 135 269 0 3
691 537
691 667
844 667
0 4 97 0 0 4096 0 0 135 270 0 3
701 520
701 676
844 676
0 0 98 0 0 4224 0 0 0 271 264 3
713 506
713 850
799 850
3 0 17 0 0 0 0 137 0 0 265 2
478 859
782 859
2 1 30 0 0 0 0 82 93 0 0 9
1396 539
1334 539
1334 667
974 667
974 904
1053 904
1053 1020
1027 1020
1027 1021
2 0 91 0 0 12416 0 130 0 0 352 7
1266 535
1239 535
1239 676
947 676
947 843
1096 843
1096 1023
2 0 92 0 0 20480 0 131 0 0 353 7
1119 539
1071 539
1071 685
934 685
934 826
1143 826
1143 1028
2 0 93 0 0 8320 0 132 0 0 350 5
981 539
919 539
919 808
1186 808
1186 1026
3 0 13 0 0 0 0 85 0 0 279 5
791 802
756 802
756 798
1236 798
1236 1023
0 0 93 0 0 0 0 0 0 280 0 2
1190 1830
1190 1998
3 9 99 0 0 4224 0 84 135 0 0 3
842 801
842 721
844 721
2 1 98 0 0 0 0 85 84 0 0 6
800 851
800 850
799 850
799 868
833 868
833 846
1 2 17 0 0 0 0 85 84 0 0 4
782 851
782 874
851 874
851 846
0 2 8 0 0 12416 0 0 79 358 0 9
1615 1127
1648 1127
1648 13
243 13
243 142
290 142
290 140
291 140
291 137
0 1 9 0 0 12416 0 0 79 354 0 7
1674 1272
1659 1272
1659 9
249 9
249 146
297 146
297 137
4 6 95 0 0 16512 0 86 130 0 0 7
635 502
635 551
680 551
680 469
1322 469
1322 535
1314 535
3 6 96 0 0 16512 0 86 131 0 0 7
641 502
641 537
691 537
691 482
1180 482
1180 539
1167 539
2 6 97 0 0 16512 0 86 132 0 0 6
647 502
647 520
701 520
701 490
1029 490
1029 539
1 6 98 0 0 0 0 86 134 0 0 7
653 502
653 506
713 506
713 499
905 499
905 527
886 527
0 0 91 0 0 0 0 0 0 273 0 2
1099 1731
1099 1997
0 0 91 0 0 0 0 0 0 274 288 2
1099 1648
1099 1731
0 0 91 0 0 0 0 0 0 327 306 2
1099 1472
1099 1648
1 4 10 0 0 12416 0 106 78 0 0 7
1652 1446
1787 1446
1787 51
346 51
346 149
312 149
312 137
0 3 11 0 0 8320 0 0 78 318 0 7
1673 1571
1793 1571
1793 46
344 46
344 146
318 146
318 137
1 2 12 0 0 8320 0 120 78 0 0 7
1673 1741
1799 1741
1799 44
342 44
342 142
324 142
324 137
1 1 13 0 0 8320 0 128 78 0 0 7
1666 1861
1805 1861
1805 40
340 40
340 138
330 138
330 137
1 1 13 0 0 0 0 128 97 0 0 4
1666 1861
1236 1861
1236 1023
1216 1023
3 0 93 0 0 0 0 124 0 0 291 3
1363 1830
1187 1830
1187 1697
2 0 92 0 0 4096 0 124 0 0 287 3
1363 1821
1143 1821
1143 1740
1 0 100 0 0 4096 0 124 0 0 360 2
1363 1812
1074 1812
4 0 101 0 0 4096 0 125 0 0 286 3
1364 1792
1167 1792
1167 1749
3 0 102 0 0 4096 0 125 0 0 305 3
1364 1783
1121 1783
1121 1657
2 0 100 0 0 4096 0 125 0 0 360 2
1364 1774
1074 1774
4 0 101 0 0 4096 0 126 0 0 308 3
1365 1749
1167 1749
1167 1610
3 0 92 0 0 4096 0 126 0 0 312 3
1365 1740
1143 1740
1143 1558
2 0 91 0 0 0 0 126 0 0 0 2
1365 1731
1096 1731
1 0 31 0 0 4096 0 126 0 0 293 3
1365 1722
1027 1722
1027 1679
4 0 33 0 0 4096 0 127 0 0 304 3
1365 1706
983 1706
983 1666
3 0 93 0 0 0 0 127 0 0 311 3
1365 1697
1187 1697
1187 1567
2 0 100 0 0 4096 0 127 0 0 360 2
1365 1688
1074 1688
1 0 31 0 0 0 0 127 0 0 313 3
1365 1679
1027 1679
1027 1549
3 0 12 0 0 0 0 121 0 0 295 2
1572 1744
1572 1743
1 3 12 0 0 0 0 120 0 0 0 3
1673 1741
1673 1743
1567 1743
0 3 93 0 0 0 0 0 124 0 0 3
1371 1831
1371 1830
1363 1830
3 1 103 0 0 4224 0 123 121 0 0 4
1481 1709
1518 1709
1518 1735
1526 1735
3 2 104 0 0 8320 0 122 121 0 0 4
1492 1793
1518 1793
1518 1753
1526 1753
5 2 105 0 0 4224 0 124 122 0 0 4
1408 1825
1438 1825
1438 1802
1446 1802
5 1 106 0 0 4224 0 125 122 0 0 4
1409 1778
1438 1778
1438 1784
1446 1784
5 2 107 0 0 4224 0 126 123 0 0 4
1410 1735
1427 1735
1427 1718
1435 1718
5 1 108 0 0 4224 0 127 123 0 0 4
1410 1692
1427 1692
1427 1700
1435 1700
3 0 92 0 0 0 0 113 0 0 326 3
1365 1524
1143 1524
1143 1481
4 0 33 0 0 0 0 116 0 0 307 3
1363 1666
983 1666
983 1619
3 0 102 0 0 0 0 116 0 0 309 3
1363 1657
1121 1657
1121 1601
2 0 91 0 0 0 0 116 0 0 0 2
1363 1648
1096 1648
4 0 33 0 0 4096 0 115 0 0 310 3
1364 1619
981 1619
981 1576
3 0 101 0 0 0 0 115 0 0 325 3
1364 1610
1167 1610
1167 1490
2 0 102 0 0 0 0 115 0 0 329 3
1364 1601
1121 1601
1121 1428
4 0 33 0 0 4096 0 114 0 0 314 3
1365 1576
981 1576
981 1533
3 0 93 0 0 0 0 114 0 0 328 3
1365 1567
1186 1567
1186 1437
2 0 92 0 0 0 0 114 0 0 303 3
1365 1558
1143 1558
1143 1524
1 0 31 0 0 0 0 114 0 0 316 3
1365 1549
1027 1549
1027 1506
4 1 33 0 0 8320 0 113 98 0 0 3
1365 1533
981 1533
981 976
2 0 100 0 0 0 0 113 0 0 360 2
1365 1515
1074 1515
1 0 31 0 0 0 0 113 0 0 334 3
1365 1506
1027 1506
1027 1366
3 0 11 0 0 0 0 119 0 0 318 2
1572 1571
1572 1571
1 3 11 0 0 0 0 112 0 0 0 3
1673 1569
1673 1571
1567 1571
3 1 109 0 0 4224 0 117 119 0 0 4
1481 1536
1518 1536
1518 1562
1526 1562
3 2 110 0 0 8320 0 118 119 0 0 4
1492 1620
1518 1620
1518 1580
1526 1580
5 2 111 0 0 4224 0 116 118 0 0 4
1408 1652
1438 1652
1438 1629
1446 1629
5 1 112 0 0 4224 0 115 118 0 0 4
1409 1605
1438 1605
1438 1611
1446 1611
5 2 113 0 0 4224 0 114 117 0 0 4
1410 1562
1427 1562
1427 1545
1435 1545
5 1 114 0 0 4224 0 113 117 0 0 4
1410 1519
1427 1519
1427 1527
1435 1527
4 0 101 0 0 4096 0 109 0 0 331 3
1367 1490
1167 1490
1167 1393
3 0 92 0 0 4096 0 109 0 0 344 3
1367 1481
1143 1481
1143 1338
2 0 91 0 0 0 0 109 0 0 333 3
1367 1472
1097 1472
1097 1375
4 0 93 0 0 0 0 110 0 0 343 3
1366 1437
1186 1437
1186 1347
3 0 102 0 0 4096 0 110 0 0 332 3
1366 1428
1121 1428
1121 1384
2 0 100 0 0 4096 0 110 0 0 360 2
1366 1419
1074 1419
4 2 101 0 0 8320 0 111 96 0 0 3
1368 1393
1167 1393
1167 1060
3 0 102 0 0 4096 0 111 0 0 346 3
1368 1384
1121 1384
1121 1302
2 0 91 0 0 0 0 111 0 0 345 3
1368 1375
1097 1375
1097 1329
1 0 31 0 0 4096 0 111 0 0 341 3
1368 1366
1027 1366
1027 1240
3 0 10 0 0 0 0 107 0 0 336 2
1551 1448
1551 1448
1 3 10 0 0 0 0 106 0 0 0 3
1652 1446
1652 1448
1546 1448
5 2 115 0 0 4224 0 109 107 0 0 4
1412 1476
1497 1476
1497 1457
1505 1457
1 3 116 0 0 8320 0 107 108 0 0 3
1505 1439
1495 1439
1495 1414
5 2 117 0 0 4224 0 110 108 0 0 2
1411 1423
1449 1423
5 1 118 0 0 4224 0 111 108 0 0 4
1413 1379
1441 1379
1441 1405
1449 1405
1 0 31 0 0 4224 0 101 0 0 342 3
1375 1240
1027 1240
1027 1204
1 2 31 0 0 0 0 104 93 0 0 3
1375 1204
1027 1204
1027 1057
3 0 93 0 0 0 0 103 0 0 350 3
1376 1347
1186 1347
1186 1222
2 0 92 0 0 4096 0 103 0 0 348 3
1376 1338
1143 1338
1143 1258
1 0 91 0 0 0 0 103 0 0 349 3
1376 1329
1097 1329
1097 1249
3 2 102 0 0 4224 0 102 95 0 0 3
1376 1302
1121 1302
1121 1060
2 0 100 0 0 4096 0 102 0 0 360 2
1376 1293
1074 1293
3 0 92 0 0 0 0 101 0 0 353 3
1375 1258
1143 1258
1143 1107
2 0 91 0 0 0 0 101 0 0 351 3
1375 1249
1096 1249
1096 1213
3 1 93 0 0 0 0 104 96 0 0 4
1375 1222
1186 1222
1186 1024
1167 1024
2 0 91 0 0 0 0 104 0 0 352 3
1375 1213
1096 1213
1096 1159
2 1 91 0 0 0 0 90 94 0 0 4
1382 1159
1096 1159
1096 1023
1074 1023
2 1 92 0 0 4224 0 92 95 0 0 4
1383 1107
1143 1107
1143 1024
1121 1024
3 1 9 0 0 0 0 87 100 0 0 3
1620 1272
1675 1272
1675 1268
3 1 119 0 0 4224 0 89 87 0 0 3
1552 1230
1552 1263
1574 1263
2 1 120 0 0 8320 0 105 89 0 0 3
1488 1222
1488 1221
1506 1221
4 0 121 0 0 0 0 104 0 0 365 2
1426 1213
1426 1213
1 3 8 0 0 0 0 99 91 0 0 3
1615 1125
1615 1127
1509 1127
0 2 32 0 0 0 0 0 97 0 0 3
1219 1058
1219 1059
1216 1059
2 0 100 0 0 4224 0 94 0 0 0 2
1074 1059
1074 1999
3 2 122 0 0 12416 0 88 87 0 0 4
1500 1317
1521 1317
1521 1281
1574 1281
4 2 123 0 0 12416 0 103 88 0 0 6
1421 1338
1419 1338
1419 1338
1446 1338
1446 1326
1454 1326
4 1 124 0 0 4224 0 102 88 0 0 4
1421 1293
1446 1293
1446 1308
1454 1308
4 2 125 0 0 12416 0 101 89 0 0 4
1420 1249
1444 1249
1444 1239
1506 1239
0 1 121 0 0 4224 0 0 105 0 0 5
1420 1213
1444 1213
1444 1221
1452 1221
1452 1222
2 3 126 0 0 4224 0 91 90 0 0 4
1463 1136
1426 1136
1426 1150
1427 1150
1 3 127 0 0 4224 0 91 92 0 0 3
1463 1118
1428 1118
1428 1098
4 4 2 0 0 128 0 131 130 0 0 3
1143 581
1290 581
1290 577
4 4 2 0 0 0 0 132 131 0 0 2
1005 581
1143 581
4 4 2 0 0 0 0 134 132 0 0 3
862 569
862 581
1005 581
1 0 2 0 0 0 0 130 0 0 372 3
1290 514
1290 411
1143 411
1 0 2 0 0 0 0 131 0 0 373 3
1143 518
1143 411
1005 411
1 0 2 0 0 0 0 132 0 0 374 3
1005 518
1005 411
864 411
1 1 2 0 0 0 0 134 129 0 0 5
862 506
862 424
864 424
864 409
826 409
4 0 94 0 0 0 0 136 0 0 376 3
793 557
796 557
796 563
0 0 94 0 0 0 0 0 0 0 380 4
797 560
796 560
796 563
797 563
3 0 94 0 0 0 0 130 0 0 378 4
1266 553
1209 553
1209 617
1105 617
3 0 94 0 0 0 0 131 0 0 379 4
1119 557
1105 557
1105 617
981 617
3 0 94 0 0 8320 0 132 0 0 380 4
981 557
981 618
797 618
797 608
1 0 94 0 0 0 0 133 0 0 381 4
820 604
820 608
797 608
797 555
0 3 94 0 0 0 0 0 134 375 0 5
793 557
793 555
797 555
797 545
838 545
8 0 128 0 0 8320 0 150 0 0 397 4
348 1016
348 1073
492 1073
492 1152
2 1 2 0 0 0 0 154 153 0 0 5
233 754
233 753
343 753
343 731
339 731
1 0 129 0 0 4096 0 1 0 0 409 2
300 841
299 841
0 1 72 0 0 0 0 0 150 386 0 3
333 917
333 953
342 953
0 0 72 0 0 0 0 0 0 389 231 4
488 919
488 917
330 917
330 919
2 2 72 0 0 0 0 139 138 0 0 4
599 908
599 919
664 919
664 912
2 0 72 0 0 0 0 140 0 0 387 3
543 907
543 919
599 919
2 0 72 0 0 0 0 137 0 0 388 3
487 904
487 919
543 919
1 0 130 0 0 12288 0 138 0 0 416 4
646 912
646 934
625 934
625 990
1 0 131 0 0 4096 0 139 0 0 415 2
581 908
581 999
1 0 132 0 0 4096 0 140 0 0 414 2
525 907
525 1008
1 0 133 0 0 4096 0 137 0 0 413 4
469 904
469 1001
470 1001
470 1016
0 0 2 0 0 0 0 0 0 395 398 3
547 1230
617 1230
617 1115
1 0 2 0 0 0 0 141 0 0 0 2
437 1230
551 1230
1 1 128 0 0 0 0 142 152 0 0 5
438 1193
552 1193
552 1192
596 1192
596 1174
1 0 128 0 0 0 0 143 0 0 396 3
439 1152
570 1152
570 1192
1 1 2 0 0 0 0 144 151 0 0 3
439 1115
640 1115
640 1129
2 0 133 0 0 8320 0 141 0 0 413 3
437 1212
531 1212
531 1016
2 0 132 0 0 8320 0 142 0 0 414 3
438 1175
503 1175
503 1007
2 0 131 0 0 8192 0 143 0 0 415 3
439 1134
478 1134
478 998
2 0 130 0 0 8192 0 144 0 0 416 3
439 1097
453 1097
453 989
1 3 134 0 0 8320 0 145 141 0 0 4
353 1171
368 1171
368 1221
382 1221
3 3 135 0 0 4224 0 145 142 0 0 3
353 1159
383 1159
383 1184
2 3 136 0 0 4224 0 145 143 0 0 3
353 1147
384 1147
384 1143
4 3 137 0 0 8320 0 145 144 0 0 4
353 1135
364 1135
364 1106
384 1106
3 5 138 0 0 8320 0 150 145 0 0 4
342 971
249 971
249 1153
302 1153
1 0 129 0 0 0 0 0 0 0 409 2
299 837
299 837
4 0 129 0 0 8320 0 150 0 0 0 3
348 980
299 980
299 834
7 0 2 0 0 0 0 150 0 0 412 2
348 1007
329 1007
6 0 2 0 0 0 0 150 0 0 412 2
348 998
329 998
1 5 2 0 0 0 0 146 150 0 0 3
329 1038
329 989
348 989
14 4 133 0 0 0 0 150 149 0 0 4
412 1016
531 1016
531 1017
631 1017
13 3 132 0 0 0 0 150 149 0 0 4
412 1007
503 1007
503 1008
631 1008
12 2 131 0 0 12416 0 150 149 0 0 4
412 998
478 998
478 999
631 999
11 1 130 0 0 12416 0 150 149 0 0 4
412 989
453 989
453 990
631 990
0 2 139 0 0 4224 0 0 150 418 0 2
135 962
348 962
3 1 139 0 0 0 0 148 147 0 0 3
84 962
135 962
135 918
33
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
46 359 297 381
55 367 287 383
29 o led aceso indica o ganhador
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
153 1426 178 1448
161 1434 169 1450
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
155 1251 214 1273
164 1259 204 1275
5 A e B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 73
794 9 808 394
797 12 804 297
73 |
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 105
33 309 810 334
39 312 803 327
105 ---------------------------------------------------------------------------------------------------------
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 105
27 0 806 25
34 3 798 18
105 ---------------------------------------------------------------------------------------------------------
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 105
36 30 813 55
42 33 806 48
105 ---------------------------------------------------------------------------------------------------------
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
442 723 525 745
451 730 515 746
8 Contador
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
388 83 417 107
398 91 406 107
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
128 15 221 39
138 23 210 39
9 Jogador 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 73
23 11 48 395
31 19 39 323
73 |
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
|
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 50
41 46 194 107
53 56 181 101
50 Clique no bot�o 
abaixo para 
sortear um valor
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
372 11 431 35
383 20 419 36
6 Placar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
712 16 789 40
722 24 778 40
7 M�quina
15 8 0 0 0 0 0 0 0 0 0 0 39
15 Liberation Sans
0 0 0 27
1010 370 1196 392
1018 374 1187 390
27 Somador 4 bits + half adder
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1541 1832 1573 1847
1553 1842 1560 1853
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1569 1713 1598 1737
1580 1721 1586 1737
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1561 1543 1592 1567
1573 1552 1579 1568
1 I
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1547 1417 1570 1441
1555 1426 1561 1442
1 H
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1562 1205 1591 1229
1573 1214 1579 1230
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1504 1094 1533 1118
1515 1103 1521 1119
1 F
15 8 0 0 0 0 0 0 0 0 0 0 39
15 Liberation Sans
0 0 0 16
85 1230 195 1251
91 1233 188 1248
16 Circuito Maquina
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
215 1364 244 1388
226 1373 232 1389
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
214 1307 243 1331
225 1316 231 1332
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
781 1649 864 1671
790 1656 854 1672
8 Contador
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
723 3082 755 3097
735 3092 742 3103
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
751 2963 780 2987
762 2971 768 2987
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
743 2793 774 2817
755 2802 761 2818
1 I
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
729 2667 752 2691
737 2676 743 2692
1 H
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
744 2455 773 2479
755 2464 761 2480
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
686 2344 715 2368
697 2353 703 2369
1 F
15 8 0 0 0 0 0 0 0 0 0 0 39
15 Liberation Sans
0 0 0 31
519 2268 687 2305
537 2279 668 2307
31 Decodificador binario 
p/ BCD
15 8 0 0 0 0 0 0 0 0 0 0 39
15 Liberation Sans
0 0 0 31
1349 1013 1517 1050
1367 1024 1498 1052
31 Decodificador binario 
p/ BCD
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
