CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1350 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
113
13 Logic Switch~
5 324 2226 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 z1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
559 0 0
2
43728.9 3
0
13 Logic Switch~
5 273 2228 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 w1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8488 0 0
2
43728.9 2
0
13 Logic Switch~
5 223 2229 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 y1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3392 0 0
2
43728.9 1
0
13 Logic Switch~
5 167 2229 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 x1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3952 0 0
2
43728.9 0
0
13 Logic Switch~
5 1081 1115 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 x3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8186 0 0
2
5.89909e-315 5.37752e-315
0
13 Logic Switch~
5 1137 1115 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 y3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6571 0 0
2
5.89909e-315 5.36716e-315
0
13 Logic Switch~
5 1187 1114 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 w3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6167 0 0
2
5.89909e-315 5.3568e-315
0
13 Logic Switch~
5 1238 1112 0 1 11
0 34
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 z3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3566 0 0
2
5.89909e-315 5.34643e-315
0
13 Logic Switch~
5 1067 1704 0 1 11
0 24
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 z2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3371 0 0
2
5.89909e-315 5.32571e-315
0
13 Logic Switch~
5 1016 1706 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 w2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4395 0 0
2
5.89909e-315 5.30499e-315
0
13 Logic Switch~
5 966 1707 0 1 11
0 39
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 y2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6822 0 0
2
5.89909e-315 5.26354e-315
0
13 Logic Switch~
5 910 1707 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 x2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8953 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 246 1459 0 1 11
0 56
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4635 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 195 1461 0 1 11
0 58
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 w
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6596 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 145 1462 0 1 11
0 54
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3813 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 89 1462 0 1 11
0 53
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 x
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5639 0 0
2
5.89909e-315 0
0
13 Logic Switch~
5 290 85 0 1 11
0 83
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
429 0 0
2
43728.9 0
0
13 Logic Switch~
5 226 83 0 1 11
0 66
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 W
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5832 0 0
2
43728.9 1
0
13 Logic Switch~
5 174 82 0 1 11
0 68
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8856 0 0
2
43728.9 2
0
13 Logic Switch~
5 116 82 0 1 11
0 71
0
0 0 21360 270
2 0V
-7 -21 7 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
469 0 0
2
43728.9 3
0
9 2-In AND~
219 1390 2269 0 3 22
0 94 95 96
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U32A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 34 0
1 U
4529 0 0
2
43728.9 0
0
9 3-In AND~
219 1641 2178 0 4 22
0 97 98 99 100
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U34A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 512 3 1 36 0
1 U
88 0 0
2
43728.9 0
0
10 2-In NAND~
219 1501 2175 0 3 22
0 101 102 103
0
0 0 624 0
6 74LS37
-14 -24 28 -16
4 U27B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 29 0
1 U
3894 0 0
2
43728.9 5
0
6 74266~
219 1412 2177 0 3 22
0 104 105 106
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 4 0
1 U
6890 0 0
2
43728.9 4
0
9 2-In AND~
219 1208 2183 0 3 22
0 107 108 109
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U21C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 23 0
1 U
3257 0 0
2
43728.9 3
0
8 2-In OR~
219 1333 2176 0 3 22
0 110 111 112
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U25A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 27 0
1 U
6612 0 0
2
43728.9 2
0
9 2-In AND~
219 1268 2181 0 3 22
0 113 114 115
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U21B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 23 0
1 U
3556 0 0
2
43728.9 1
0
9 2-In XOR~
219 1561 2176 0 3 22
0 116 117 118
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U29A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 31 0
1 U
9143 0 0
2
43728.9 0
0
4 LED~
171 628 2474 0 2 2
10 3 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8186 0 0
2
43728.9 1
0
7 Ground~
168 628 2506 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3754 0 0
2
43728.9 0
0
8 2-In OR~
219 564 2448 0 3 22
0 5 4 3
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U30A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
8708 0 0
2
43728.9 0
0
8 2-In OR~
219 472 2385 0 3 22
0 7 6 5
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U25D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
3338 0 0
2
43728.9 0
0
9 2-In AND~
219 464 2509 0 3 22
0 9 8 4
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U28C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
5546 0 0
2
43728.9 0
0
10 2-In NAND~
219 390 2491 0 3 22
0 10 11 9
0
0 0 624 0
6 74LS37
-14 -24 28 -16
4 U27C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 29 0
1 U
3295 0 0
2
43728.9 0
0
9 2-In AND~
219 388 2423 0 3 22
0 13 12 6
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U28B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
4923 0 0
2
43728.9 0
0
9 2-In XOR~
219 380 2358 0 3 22
0 15 14 7
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U29B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
3248 0 0
2
43728.9 0
0
9 Inverter~
13 253 2292 0 2 22
0 10 13
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U24E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 26 0
1 U
3139 0 0
2
43728.9 7
0
9 Inverter~
13 303 2293 0 2 22
0 12 11
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U24D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 26 0
1 U
3285 0 0
2
43728.9 6
0
9 Inverter~
13 137 2286 0 2 22
0 15 8
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U24C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 26 0
1 U
336 0 0
2
43728.9 5
0
9 Inverter~
13 202 2287 0 2 22
0 14 16
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U24B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 26 0
1 U
6582 0 0
2
43728.9 4
0
4 LED~
171 1437 1991 0 2 2
10 17 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3546 0 0
2
43728.9 1
0
7 Ground~
168 1437 2023 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
893 0 0
2
43728.9 0
0
8 2-In OR~
219 1367 1952 0 3 22
0 18 19 17
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U25C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
8998 0 0
2
43728.9 0
0
8 2-In OR~
219 1289 1864 0 3 22
0 21 20 18
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U25B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 27 0
1 U
5979 0 0
2
43728.9 0
0
9 2-In AND~
219 1202 2035 0 3 22
0 23 22 19
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U28A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
3835 0 0
2
43728.9 0
0
10 2-In NAND~
219 1135 1992 0 3 22
0 25 24 23
0
0 0 624 0
6 74LS37
-14 -24 28 -16
4 U27A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
750 0 0
2
43728.9 0
0
9 2-In AND~
219 1215 1918 0 3 22
0 27 26 20
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U21D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 23 0
1 U
849 0 0
2
43728.9 0
0
6 74266~
219 1125 1881 0 3 22
0 28 24 27
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4693 0 0
2
43728.9 0
0
9 3-In AND~
219 1129 1818 0 4 22
0 25 29 24 21
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U26A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 28 0
1 U
4775 0 0
2
43728.9 0
0
9 Inverter~
13 1116 1173 0 2 22
0 36 31
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U24A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 26 0
1 U
9572 0 0
2
5.89909e-315 5.32571e-315
0
9 Inverter~
13 1051 1172 0 2 22
0 37 30
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U23F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 25 0
1 U
3761 0 0
2
5.89909e-315 5.30499e-315
0
9 Inverter~
13 1217 1179 0 2 22
0 34 33
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U23E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 25 0
1 U
6765 0 0
2
5.89909e-315 5.26354e-315
0
9 Inverter~
13 1167 1178 0 2 22
0 35 32
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U23D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 25 0
1 U
7938 0 0
2
5.89909e-315 0
0
9 Inverter~
13 996 1770 0 2 22
0 28 29
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U23C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 25 0
1 U
55 0 0
2
5.89909e-315 5.37752e-315
0
9 Inverter~
13 1046 1771 0 2 22
0 24 38
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U23B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 25 0
1 U
5610 0 0
2
5.89909e-315 5.36716e-315
0
9 Inverter~
13 880 1764 0 2 22
0 25 26
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U23A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 25 0
1 U
3322 0 0
2
5.89909e-315 5.3568e-315
0
9 Inverter~
13 945 1765 0 2 22
0 39 22
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U20F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 22 0
1 U
5914 0 0
2
5.89909e-315 5.34643e-315
0
4 LED~
171 942 1481 0 2 2
10 119 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 512 1 0 0 0
1 D
8748 0 0
2
5.89909e-315 5.26354e-315
0
7 Ground~
168 942 1513 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5830 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 610 1711 0 3 22
0 41 42 40
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U22D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 24 0
1 U
9153 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 520 1632 0 3 22
0 44 43 41
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U22B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 24 0
1 U
9220 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 444 1821 0 3 22
0 46 45 42
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U22A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
7901 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 436 1701 0 3 22
0 48 47 43
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
4571 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 427 1583 0 3 22
0 50 49 44
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
7796 0 0
2
5.89909e-315 0
0
9 3-In AND~
219 320 1847 0 4 22
0 53 52 51 45
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 18 0
1 U
3907 0 0
2
5.89909e-315 0
0
9 3-In AND~
219 321 1793 0 4 22
0 56 55 54 46
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 18 0
1 U
4389 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 324 1729 0 3 22
0 57 52 47
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 23 0
1 U
7762 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 324 1671 0 3 22
0 53 57 48
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
6723 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 324 1615 0 3 22
0 54 58 49
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6871 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 322 1553 0 3 22
0 55 58 50
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
4198 0 0
2
5.89909e-315 0
0
9 Inverter~
13 175 1525 0 2 22
0 58 51
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U20A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 22 0
1 U
970 0 0
2
5.89909e-315 0
0
9 Inverter~
13 225 1526 0 2 22
0 56 57
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
319 0 0
2
5.89909e-315 0
0
9 Inverter~
13 59 1519 0 2 22
0 53 55
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
3663 0 0
2
5.89909e-315 0
0
9 Inverter~
13 124 1520 0 2 22
0 54 52
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
3512 0 0
2
5.89909e-315 0
0
7 Ground~
168 680 1796 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7555 0 0
2
5.89909e-315 0
0
4 LED~
171 680 1764 0 2 2
10 40 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9776 0 0
2
5.89909e-315 0
0
9 3-In AND~
219 405 1322 0 4 22
0 120 121 122 123
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 512 3 1 18 0
1 U
6596 0 0
2
5.89909e-315 0
0
9 2-In AND~
219 343 1324 0 3 22
0 124 125 126
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 5 0
1 U
6750 0 0
2
5.89909e-315 0
0
9 Inverter~
13 274 1323 0 2 22
0 127 128
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U10C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 3 12 0
1 U
9636 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 196 1324 0 3 22
0 129 130 131
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 15 0
1 U
5369 0 0
2
5.89909e-315 0
0
7 Ground~
168 674 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8555 0 0
2
5.89909e-315 0
0
9 CC 7-Seg~
183 607 384 0 17 19
10 65 64 63 62 61 60 59 132 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4690 0 0
2
5.89909e-315 5.26354e-315
0
8 2-In OR~
219 515 1013 0 3 22
0 71 73 76
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
9145 0 0
2
5.89909e-315 5.30499e-315
0
8 2-In OR~
219 508 1124 0 3 22
0 75 74 72
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
5246 0 0
2
5.89909e-315 5.32571e-315
0
8 2-In OR~
219 579 1073 0 3 22
0 76 72 59
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
9111 0 0
2
5.89909e-315 5.34643e-315
0
9 2-In AND~
219 416 1034 0 3 22
0 66 67 73
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
6717 0 0
2
5.89909e-315 5.3568e-315
0
9 2-In AND~
219 416 1092 0 3 22
0 68 69 75
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
3487 0 0
2
5.89909e-315 5.36716e-315
0
9 2-In AND~
219 415 1151 0 3 22
0 66 70 74
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
9604 0 0
2
5.89909e-315 5.37752e-315
0
8 2-In OR~
219 557 892 0 3 22
0 78 77 60
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3921 0 0
2
5.89909e-315 5.38788e-315
0
8 2-In OR~
219 482 930 0 3 22
0 80 79 77
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
8146 0 0
2
5.89909e-315 5.39306e-315
0
8 2-In OR~
219 485 855 0 3 22
0 81 71 78
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
4506 0 0
2
5.89909e-315 5.39824e-315
0
9 2-In AND~
219 409 832 0 3 22
0 68 70 81
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
5386 0 0
2
5.89909e-315 5.40342e-315
0
9 2-In AND~
219 408 899 0 3 22
0 68 69 80
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
7847 0 0
2
5.89909e-315 5.4086e-315
0
9 2-In AND~
219 405 958 0 3 22
0 69 70 79
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
9261 0 0
2
5.89909e-315 5.41378e-315
0
9 2-In AND~
219 553 746 0 3 22
0 82 70 61
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
8231 0 0
2
5.89909e-315 5.41896e-315
0
8 2-In OR~
219 446 717 0 3 22
0 67 66 82
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3756 0 0
2
5.89909e-315 5.42414e-315
0
9 3-In AND~
219 399 636 0 4 22
0 69 83 68 86
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 6 0
1 U
6760 0 0
2
43728.9 4
0
8 3-In OR~
219 556 553 0 4 22
0 88 87 86 62
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
351 0 0
2
43728.9 5
0
8 3-In OR~
219 485 470 0 4 22
0 71 85 84 88
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
5352 0 0
2
43728.9 6
0
9 2-In AND~
219 403 481 0 3 22
0 70 66 85
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
485 0 0
2
43728.9 7
0
9 2-In AND~
219 402 530 0 3 22
0 67 70 84
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
452 0 0
2
43728.9 8
0
9 2-In AND~
219 397 588 0 3 22
0 67 66 87
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
643 0 0
2
43728.9 9
0
8 2-In OR~
219 495 385 0 3 22
0 68 89 63
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
5563 0 0
2
43728.9 10
0
8 2-In OR~
219 412 411 0 3 22
0 69 83 89
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
934 0 0
2
43728.9 11
0
6 74266~
219 369 352 0 3 22
0 66 83 90
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3240 0 0
2
43728.9 12
0
8 2-In OR~
219 491 303 0 3 22
0 67 90 64
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3233 0 0
2
43728.9 13
0
8 2-In OR~
219 388 188 0 3 22
0 71 66 92
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3635 0 0
2
43728.9 14
0
8 2-In OR~
219 485 221 0 3 22
0 92 91 65
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3547 0 0
2
43728.9 15
0
6 74266~
219 390 264 0 3 22
0 68 83 91
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
483 0 0
2
43728.9 16
0
9 Inverter~
13 260 136 0 2 22
0 83 70
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
6126 0 0
2
43728.9 17
0
9 Inverter~
13 199 134 0 2 22
0 66 69
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
7368 0 0
2
43728.9 18
0
9 Inverter~
13 143 131 0 2 22
0 68 67
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3925 0 0
2
43728.9 19
0
9 Inverter~
13 82 132 0 2 22
0 71 93
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
6187 0 0
2
43728.9 20
0
184
3 1 3 0 0 4224 0 31 29 0 0 3
597 2448
628 2448
628 2464
1 2 2 0 0 4096 0 30 29 0 0 2
628 2500
628 2484
3 2 4 0 0 4224 0 33 31 0 0 4
485 2509
543 2509
543 2457
551 2457
3 1 5 0 0 8320 0 32 31 0 0 4
505 2385
543 2385
543 2439
551 2439
3 2 6 0 0 4224 0 35 32 0 0 4
409 2423
451 2423
451 2394
459 2394
3 1 7 0 0 4224 0 36 32 0 0 4
413 2358
451 2358
451 2376
459 2376
2 0 8 0 0 4096 0 33 0 0 15 2
440 2518
140 2518
3 1 9 0 0 4224 0 34 33 0 0 4
417 2491
432 2491
432 2500
440 2500
1 0 10 0 0 4096 0 34 0 0 24 2
366 2482
273 2482
2 0 11 0 0 4096 0 34 0 0 18 2
366 2500
306 2500
2 0 12 0 0 4096 0 35 0 0 23 2
364 2432
324 2432
1 0 13 0 0 4096 0 35 0 0 17 2
364 2414
256 2414
2 0 14 0 0 4096 0 36 0 0 25 2
364 2367
223 2367
1 0 15 0 0 4096 0 36 0 0 26 2
364 2349
167 2349
2 0 8 0 0 4224 0 39 0 0 0 2
140 2304
140 2703
2 0 16 0 0 4224 0 40 0 0 0 2
205 2305
205 2703
2 0 13 0 0 4224 0 37 0 0 0 2
256 2310
256 2702
2 0 11 0 0 4224 0 38 0 0 0 2
306 2311
306 2702
1 0 12 0 0 0 0 38 0 0 23 3
306 2275
306 2250
324 2250
1 0 10 0 0 0 0 37 0 0 24 3
256 2274
256 2250
273 2250
1 0 14 0 0 0 0 40 0 0 25 3
205 2269
205 2251
223 2251
1 0 15 0 0 0 0 39 0 0 26 3
140 2268
140 2253
167 2253
1 0 12 0 0 4224 0 1 0 0 0 2
324 2238
324 2701
1 0 10 0 0 4224 0 2 0 0 0 2
273 2240
273 2701
1 0 14 0 0 4224 0 3 0 0 0 2
223 2241
223 2704
1 0 15 0 0 4224 0 4 0 0 0 2
167 2241
167 2702
3 1 17 0 0 4224 0 43 41 0 0 3
1400 1952
1437 1952
1437 1981
1 2 2 0 0 0 0 42 41 0 0 2
1437 2017
1437 2001
3 1 18 0 0 8320 0 44 43 0 0 4
1322 1864
1349 1864
1349 1943
1354 1943
3 2 19 0 0 4224 0 45 43 0 0 4
1223 2035
1349 2035
1349 1961
1354 1961
3 2 20 0 0 8320 0 47 44 0 0 4
1236 1918
1262 1918
1262 1873
1276 1873
4 1 21 0 0 4224 0 49 44 0 0 4
1150 1818
1262 1818
1262 1855
1276 1855
2 0 22 0 0 4096 0 45 0 0 57 2
1178 2044
948 2044
3 1 23 0 0 8320 0 46 45 0 0 4
1162 1992
1170 1992
1170 2026
1178 2026
2 0 24 0 0 4096 0 46 0 0 64 2
1111 2001
1067 2001
1 0 25 0 0 4096 0 46 0 0 67 2
1111 1983
910 1983
2 0 26 0 0 4096 0 47 0 0 56 2
1191 1927
883 1927
3 1 27 0 0 8320 0 48 47 0 0 4
1164 1881
1183 1881
1183 1909
1191 1909
2 0 24 0 0 0 0 48 0 0 64 2
1109 1890
1067 1890
1 0 28 0 0 4096 0 48 0 0 65 2
1109 1872
1016 1872
3 0 24 0 0 0 0 49 0 0 64 2
1105 1827
1067 1827
2 0 29 0 0 4096 0 49 0 0 58 2
1105 1818
999 1818
1 0 25 0 0 0 0 49 0 0 67 2
1105 1809
910 1809
2 0 30 0 0 4224 0 51 0 0 0 2
1054 1190
1054 1589
2 0 31 0 0 4224 0 50 0 0 0 2
1119 1191
1119 1589
2 0 32 0 0 4224 0 53 0 0 0 2
1170 1196
1170 1588
2 0 33 0 0 4224 0 52 0 0 0 2
1220 1197
1220 1588
1 0 34 0 0 4096 0 52 0 0 52 3
1220 1161
1220 1136
1238 1136
1 0 35 0 0 4096 0 53 0 0 53 3
1170 1160
1170 1136
1187 1136
1 0 36 0 0 4096 0 50 0 0 54 3
1119 1155
1119 1137
1137 1137
1 0 37 0 0 8192 0 51 0 0 55 3
1054 1154
1054 1139
1081 1139
1 0 34 0 0 4224 0 8 0 0 0 2
1238 1124
1238 1587
1 0 35 0 0 4224 0 7 0 0 0 2
1187 1126
1187 1587
1 0 36 0 0 4224 0 6 0 0 0 2
1137 1127
1137 1590
1 0 37 0 0 4224 0 5 0 0 0 2
1081 1127
1081 1588
2 0 26 0 0 4224 0 56 0 0 0 2
883 1782
883 2181
2 0 22 0 0 4224 0 57 0 0 0 2
948 1783
948 2181
2 0 29 0 0 4224 0 54 0 0 0 2
999 1788
999 2180
2 0 38 0 0 4224 0 55 0 0 0 2
1049 1789
1049 2180
1 0 24 0 0 0 0 55 0 0 64 3
1049 1753
1049 1728
1067 1728
1 0 28 0 0 0 0 54 0 0 65 3
999 1752
999 1728
1016 1728
1 0 39 0 0 4096 0 57 0 0 66 3
948 1747
948 1729
966 1729
1 0 25 0 0 0 0 56 0 0 67 3
883 1746
883 1731
910 1731
1 0 24 0 0 4224 0 9 0 0 0 2
1067 1716
1067 2179
1 0 28 0 0 4224 0 10 0 0 0 2
1016 1718
1016 2179
1 0 39 0 0 4224 0 11 0 0 0 2
966 1719
966 2182
1 0 25 0 0 4224 0 12 0 0 0 2
910 1719
910 2180
3 1 40 0 0 8320 0 60 76 0 0 3
643 1711
680 1711
680 1754
1 2 2 0 0 0 0 59 58 0 0 2
942 1507
942 1491
1 2 2 0 0 0 0 75 76 0 0 2
680 1790
680 1774
3 1 41 0 0 8320 0 61 60 0 0 4
553 1632
589 1632
589 1702
597 1702
3 2 42 0 0 8320 0 62 60 0 0 4
477 1821
563 1821
563 1720
597 1720
3 2 43 0 0 8320 0 63 61 0 0 4
469 1701
499 1701
499 1641
507 1641
3 1 44 0 0 8320 0 64 61 0 0 4
460 1583
499 1583
499 1623
507 1623
4 2 45 0 0 4224 0 65 62 0 0 4
341 1847
423 1847
423 1830
431 1830
4 1 46 0 0 4224 0 66 62 0 0 4
342 1793
423 1793
423 1812
431 1812
3 2 47 0 0 4224 0 67 63 0 0 4
345 1729
417 1729
417 1710
423 1710
3 1 48 0 0 4224 0 68 63 0 0 4
345 1671
417 1671
417 1692
423 1692
3 2 49 0 0 4224 0 69 64 0 0 4
345 1615
407 1615
407 1592
414 1592
3 1 50 0 0 4224 0 70 64 0 0 4
343 1553
407 1553
407 1574
414 1574
3 0 51 0 0 4096 0 65 0 0 97 2
296 1856
178 1856
2 0 52 0 0 4096 0 65 0 0 96 2
296 1847
127 1847
1 0 53 0 0 4096 0 68 0 0 106 2
300 1662
89 1662
1 0 53 0 0 0 0 65 0 0 106 2
296 1838
89 1838
3 0 54 0 0 4096 0 66 0 0 105 2
297 1802
145 1802
2 0 55 0 0 4096 0 66 0 0 95 2
297 1793
62 1793
1 0 56 0 0 4096 0 66 0 0 103 2
297 1784
246 1784
2 0 52 0 0 4096 0 67 0 0 96 2
300 1738
127 1738
1 0 57 0 0 4096 0 67 0 0 98 2
300 1720
228 1720
2 0 57 0 0 0 0 68 0 0 98 2
300 1680
228 1680
2 0 58 0 0 4096 0 69 0 0 104 2
300 1624
195 1624
1 0 54 0 0 4096 0 69 0 0 105 2
300 1606
145 1606
2 0 58 0 0 0 0 70 0 0 104 2
298 1562
195 1562
0 1 55 0 0 8192 0 0 70 95 0 3
62 1543
62 1544
298 1544
2 0 55 0 0 4224 0 73 0 0 0 2
62 1537
62 1888
2 0 52 0 0 4224 0 74 0 0 0 2
127 1538
127 1889
2 0 51 0 0 4224 0 71 0 0 0 2
178 1543
178 1894
2 0 57 0 0 4224 0 72 0 0 0 2
228 1544
228 1893
1 0 56 0 0 0 0 72 0 0 103 3
228 1508
228 1483
246 1483
1 0 58 0 0 0 0 71 0 0 104 3
178 1507
178 1483
195 1483
1 0 54 0 0 0 0 74 0 0 105 3
127 1502
127 1484
145 1484
1 0 53 0 0 0 0 73 0 0 106 3
62 1501
62 1486
89 1486
1 0 56 0 0 4224 0 13 0 0 0 2
246 1471
246 1894
1 0 58 0 0 4224 0 14 0 0 0 2
195 1473
195 1891
1 0 54 0 0 4224 0 15 0 0 0 2
145 1474
145 1890
1 0 53 0 0 4224 0 16 0 0 0 2
89 1474
89 1890
7 3 59 0 0 4224 0 82 85 0 0 3
622 420
622 1073
612 1073
6 3 60 0 0 4224 0 82 89 0 0 3
616 420
616 892
590 892
5 3 61 0 0 4224 0 82 95 0 0 3
610 420
610 746
574 746
4 4 62 0 0 4224 0 82 98 0 0 3
604 420
604 553
589 553
3 3 63 0 0 8320 0 82 103 0 0 5
598 420
598 430
541 430
541 385
528 385
2 3 64 0 0 12416 0 82 106 0 0 5
592 420
592 425
537 425
537 303
524 303
1 3 65 0 0 8320 0 82 108 0 0 4
586 420
533 420
533 221
518 221
1 9 2 0 0 4224 0 81 82 0 0 4
674 426
674 330
607 330
607 342
1 0 66 0 0 4096 0 86 0 0 177 2
392 1025
226 1025
2 0 67 0 0 4096 0 86 0 0 180 2
392 1043
146 1043
1 0 68 0 0 4096 0 87 0 0 181 2
392 1083
174 1083
2 0 69 0 0 4096 0 87 0 0 176 2
392 1101
202 1101
2 0 70 0 0 4096 0 88 0 0 174 2
391 1160
263 1160
1 0 66 0 0 0 0 88 0 0 177 2
391 1142
226 1142
1 0 71 0 0 4096 0 83 0 0 184 2
502 1004
116 1004
3 2 72 0 0 8320 0 84 85 0 0 4
541 1124
558 1124
558 1082
566 1082
3 2 73 0 0 4224 0 86 83 0 0 4
437 1034
471 1034
471 1022
502 1022
3 2 74 0 0 4224 0 88 84 0 0 4
436 1151
476 1151
476 1133
495 1133
3 1 75 0 0 4224 0 87 84 0 0 4
437 1092
476 1092
476 1115
495 1115
3 1 76 0 0 4224 0 83 85 0 0 3
548 1013
548 1064
566 1064
2 0 70 0 0 0 0 94 0 0 174 2
381 967
263 967
2 0 69 0 0 0 0 93 0 0 176 2
384 908
202 908
1 0 69 0 0 0 0 94 0 0 176 2
381 949
202 949
2 0 70 0 0 0 0 92 0 0 174 2
385 841
263 841
1 0 68 0 0 0 0 92 0 0 181 2
385 823
174 823
2 0 71 0 0 0 0 91 0 0 184 2
472 864
116 864
3 2 77 0 0 8320 0 90 89 0 0 4
515 930
536 930
536 901
544 901
3 1 78 0 0 8320 0 91 89 0 0 4
518 855
536 855
536 883
544 883
3 2 79 0 0 4224 0 94 90 0 0 4
426 958
461 958
461 939
469 939
3 1 80 0 0 4224 0 93 90 0 0 4
429 899
461 899
461 921
469 921
3 1 81 0 0 8320 0 92 91 0 0 3
430 832
430 846
472 846
0 1 68 0 0 0 0 0 93 181 0 2
174 890
384 890
0 2 70 0 0 4096 0 0 95 174 0 4
263 781
513 781
513 755
529 755
3 1 82 0 0 4224 0 96 95 0 0 4
479 717
512 717
512 737
529 737
0 2 66 0 0 4096 0 0 96 177 0 4
226 741
396 741
396 726
433 726
0 1 67 0 0 4096 0 0 96 180 0 4
146 693
396 693
396 708
433 708
3 0 68 0 0 0 0 97 0 0 181 2
375 645
174 645
2 0 83 0 0 4096 0 97 0 0 173 2
375 636
290 636
1 0 69 0 0 0 0 97 0 0 176 2
375 627
202 627
2 0 66 0 0 0 0 102 0 0 177 2
373 597
226 597
1 0 67 0 0 0 0 102 0 0 180 2
373 579
146 579
2 0 70 0 0 0 0 101 0 0 174 2
378 539
263 539
1 0 70 0 0 0 0 100 0 0 174 2
379 472
263 472
1 0 67 0 0 0 0 101 0 0 180 2
378 521
146 521
2 0 66 0 0 0 0 100 0 0 177 2
379 490
226 490
3 3 84 0 0 8320 0 101 99 0 0 4
423 530
452 530
452 479
472 479
3 2 85 0 0 12416 0 100 99 0 0 4
424 481
440 481
440 470
473 470
1 0 71 0 0 0 0 99 0 0 184 2
472 461
116 461
4 3 86 0 0 4224 0 97 98 0 0 4
420 636
520 636
520 562
543 562
3 2 87 0 0 4224 0 102 98 0 0 4
418 588
495 588
495 553
544 553
4 1 88 0 0 8320 0 99 98 0 0 4
518 470
535 470
535 544
543 544
1 0 69 0 0 4096 0 104 0 0 176 2
399 402
202 402
2 0 83 0 0 4096 0 104 0 0 173 2
399 420
290 420
1 0 68 0 0 4096 0 103 0 0 181 2
482 376
174 376
3 2 89 0 0 4224 0 104 103 0 0 4
445 411
474 411
474 394
482 394
2 0 83 0 0 0 0 105 0 0 173 2
353 361
290 361
1 0 66 0 0 0 0 105 0 0 177 2
353 343
226 343
1 0 67 0 0 4096 0 106 0 0 180 2
478 294
146 294
3 2 90 0 0 8320 0 105 106 0 0 3
408 352
408 312
478 312
2 0 83 0 0 0 0 109 0 0 173 2
374 273
290 273
1 0 71 0 0 0 0 107 0 0 184 2
375 179
116 179
3 2 91 0 0 4224 0 109 108 0 0 4
429 264
464 264
464 230
472 230
0 1 68 0 0 0 0 0 109 181 0 4
174 220
367 220
367 255
374 255
0 2 66 0 0 0 0 0 107 177 0 4
226 260
349 260
349 197
375 197
3 1 92 0 0 4224 0 107 108 0 0 4
421 188
452 188
452 212
472 212
0 1 83 0 0 0 0 0 110 173 0 3
290 109
263 109
263 118
1 0 83 0 0 4224 0 17 0 0 0 2
290 97
290 1209
2 0 70 0 0 4224 0 110 0 0 0 2
263 154
263 1212
1 0 66 0 0 0 0 111 0 0 177 2
202 116
226 116
2 0 69 0 0 4224 0 111 0 0 0 2
202 152
202 1215
1 0 66 0 0 4224 0 18 0 0 0 2
226 95
226 1212
1 0 68 0 0 0 0 112 0 0 181 2
146 113
174 113
1 0 71 0 0 0 0 113 0 0 184 2
85 114
116 114
2 0 67 0 0 4224 0 112 0 0 0 2
146 149
146 1215
1 0 68 0 0 4224 0 19 0 0 0 2
174 94
174 1214
1 0 68 0 0 0 0 19 0 0 0 2
174 94
174 656
2 0 93 0 0 4224 0 113 0 0 0 2
85 150
85 1217
1 0 71 0 0 4224 0 20 0 0 0 2
116 94
116 1216
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
398 2274 659 2298
408 2282 648 2298
30 C = X'(WZ')' + W'Z + (X XOR Y)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
391 2244 420 2268
401 2252 409 2268
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
290 2193 319 2217
300 2201 308 2217
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 35
888 1634 1189 1658
898 1642 1178 1658
35 b = XW'Z + X'( W NXOR Z) + Y' (XY)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 499 610 523
593 507 601 523
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
518 350 547 374
528 358 536 374
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
529 269 554 293
537 277 545 293
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
527 187 556 211
537 195 545 211
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1204 1079 1233 1103
1214 1087 1222 1103
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1299 676 1376 700
1309 684 1365 700
7 SAIDA D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
576 691 605 715
586 699 594 715
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
581 844 610 868
591 852 599 868
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 1006 614 1030
595 1014 603 1030
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
47 1298 116 1322
57 1306 105 1322
6 a hexa
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
71 1366 412 1390
81 1374 401 1390
40 a = x'w + yw + xz' + z'y' + zx'y + xy'w'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
901 1605 978 1629
911 1613 967 1629
7 saida b
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
