CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 2 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
25
7 Ground~
168 761 90 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
43785.6 0
0
7 Ground~
168 20 192 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
391 0 0
2
43785.6 0
0
7 Pulser~
4 63 170 0 10 12
0 2 2 4 26 0 0 5 5 4
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3124 0 0
2
43785.6 0
0
7 Ground~
168 261 29 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3421 0 0
2
43785.6 0
0
5 4013~
219 378 146 0 6 22
0 2 6 7 5 6 9
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 8 0
1 U
8157 0 0
2
43785.6 0
0
5 4013~
219 261 147 0 6 22
0 2 7 8 5 7 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 2 7 0
1 U
5572 0 0
2
43785.6 0
0
5 4013~
219 119 146 0 6 22
0 2 8 4 5 8 10
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 0 2 1 7 0
1 U
8901 0 0
2
43785.6 0
0
7 Ground~
168 57 402 0 1 3
0 2
0
0 0 53360 602
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
5.89916e-315 0
0
2 +V
167 29 365 0 1 3
0 11
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4747 0 0
2
5.89916e-315 0
0
6 74LS85
106 276 389 0 14 29
0 2 9 3 10 2 11 11 11 27
28 29 30 5 31
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U7
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
972 0 0
2
5.89916e-315 0
0
2 +V
167 587 309 0 1 3
0 12
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.89916e-315 0
0
5 4049~
219 481 575 0 2 22
0 10 15
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6C
-12 14 9 22
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 6 0
1 U
9998 0 0
2
5.89916e-315 0
0
5 4049~
219 481 502 0 2 22
0 9 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 6 0
1 U
3536 0 0
2
5.89916e-315 0
0
5 4049~
219 483 547 0 2 22
0 3 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 6 0
1 U
4597 0 0
2
5.89916e-315 0
0
5 4081~
219 639 421 0 3 22
0 10 13 25
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3835 0 0
2
5.89916e-315 5.39306e-315
0
5 4081~
219 637 467 0 3 22
0 3 15 24
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
3670 0 0
2
5.89916e-315 5.38788e-315
0
5 4081~
219 636 511 0 3 22
0 13 15 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
5616 0 0
2
5.89916e-315 5.37752e-315
0
5 4081~
219 636 661 0 3 22
0 9 13 20
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
9323 0 0
2
5.89916e-315 5.36716e-315
0
5 4081~
219 640 614 0 3 22
0 14 10 21
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
317 0 0
2
5.89916e-315 5.3568e-315
0
5 4081~
219 639 571 0 3 22
0 3 9 22
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3108 0 0
2
5.89916e-315 5.34643e-315
0
5 4071~
219 776 421 0 3 22
0 3 25 19
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
5.89916e-315 5.32571e-315
0
5 4071~
219 779 464 0 3 22
0 25 24 18
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
5.89916e-315 5.30499e-315
0
5 4071~
219 787 564 0 3 22
0 21 20 16
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
7876 0 0
2
5.89916e-315 5.26354e-315
0
5 4071~
219 784 521 0 3 22
0 23 22 17
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
6369 0 0
2
5.89916e-315 0
0
9 CC 7-Seg~
183 844 129 0 17 19
10 12 19 18 17 12 12 16 32 2
1 1 0 0 1 1 1 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9172 0 0
2
5.89916e-315 0
0
54
0 0 3 0 0 16384 0 0 0 18 40 6
303 111
321 111
321 268
411 268
411 547
433 547
1 9 2 0 0 8192 0 1 25 0 0 4
761 84
761 54
844 54
844 87
3 3 4 0 0 4224 0 3 7 0 0 3
87 161
87 128
95 128
1 0 2 0 0 0 0 2 0 0 5 3
20 186
20 165
33 165
1 2 2 0 0 0 0 3 3 0 0 3
39 161
33 161
33 170
0 4 5 0 0 4096 0 0 7 7 0 3
263 203
119 203
119 152
0 4 5 0 0 0 0 0 6 8 0 3
378 203
261 203
261 153
13 4 5 0 0 8320 0 10 5 0 0 3
308 416
378 416
378 152
2 5 6 0 0 12416 0 5 5 0 0 6
354 110
342 110
342 76
447 76
447 128
408 128
2 0 7 0 0 12416 0 6 0 0 15 5
237 111
219 111
219 73
332 73
332 129
2 0 8 0 0 12416 0 7 0 0 16 5
95 110
82 110
82 72
196 72
196 129
1 0 2 0 0 0 0 6 0 0 13 2
261 90
261 49
0 1 2 0 0 4096 0 0 5 14 0 3
261 49
378 49
378 89
1 1 2 0 0 8192 0 7 4 0 0 4
119 89
119 49
261 49
261 37
5 3 7 0 0 0 0 6 5 0 0 4
291 129
339 129
339 128
354 128
5 3 8 0 0 0 0 7 6 0 0 4
149 128
164 128
164 129
237 129
6 2 9 0 0 12416 0 5 10 0 0 6
402 110
429 110
429 305
160 305
160 371
244 371
6 3 3 0 0 128 0 6 10 0 0 6
285 111
303 111
303 324
212 324
212 380
244 380
6 4 10 0 0 8192 0 7 10 0 0 4
143 110
182 110
182 389
244 389
1 0 2 0 0 0 0 10 0 0 21 3
244 362
119 362
119 398
1 5 2 0 0 12416 0 8 10 0 0 4
64 403
79 403
79 398
244 398
0 1 11 0 0 4096 0 0 9 23 0 3
122 423
29 423
29 374
0 7 11 0 0 8320 0 0 10 24 0 3
122 423
122 416
244 416
6 8 11 0 0 0 0 10 10 0 0 4
244 407
122 407
122 425
244 425
1 0 12 0 0 8320 0 11 0 0 54 5
587 318
587 369
807 369
807 176
823 176
0 2 13 0 0 4224 0 0 18 33 0 3
539 547
539 670
612 670
0 1 9 0 0 0 0 0 18 31 0 3
559 605
559 652
612 652
1 2 14 0 0 8320 0 19 13 0 0 6
616 605
601 605
601 511
547 511
547 502
502 502
0 2 10 0 0 128 0 0 19 39 0 3
449 575
449 623
616 623
0 1 3 0 0 0 0 0 20 38 0 3
585 396
585 562
615 562
0 2 9 0 0 128 0 0 20 41 0 5
438 502
438 605
589 605
589 580
615 580
0 2 15 0 0 8192 0 0 17 34 0 4
530 575
574 575
574 520
612 520
0 1 13 0 0 0 0 0 17 37 0 4
513 547
563 547
563 502
612 502
2 2 15 0 0 8320 0 12 16 0 0 4
502 575
530 575
530 476
613 476
1 0 3 0 0 0 0 16 0 0 38 2
613 458
446 458
0 1 10 0 0 0 0 0 15 39 0 3
457 575
457 412
615 412
2 2 13 0 0 0 0 14 15 0 0 4
504 547
513 547
513 430
615 430
0 1 3 0 0 8320 0 0 21 40 0 5
446 547
446 396
730 396
730 412
763 412
0 1 10 0 0 4224 0 0 12 19 0 3
174 110
174 575
466 575
0 1 3 0 0 0 0 0 14 0 0 2
430 547
468 547
0 1 9 0 0 0 0 0 13 17 0 6
427 110
451 110
451 364
428 364
428 502
466 502
3 7 16 0 0 8320 0 23 25 0 0 3
820 564
859 564
859 165
4 3 17 0 0 4224 0 25 24 0 0 3
841 165
841 521
817 521
3 3 18 0 0 8320 0 22 25 0 0 3
812 464
835 464
835 165
3 2 19 0 0 8320 0 21 25 0 0 3
809 421
829 421
829 165
2 3 20 0 0 8320 0 23 18 0 0 4
774 573
709 573
709 661
657 661
1 3 21 0 0 4224 0 23 19 0 0 4
774 555
699 555
699 614
661 614
2 3 22 0 0 4224 0 24 20 0 0 4
771 530
678 530
678 571
660 571
3 1 23 0 0 8320 0 17 24 0 0 3
657 511
657 512
771 512
3 2 24 0 0 4224 0 16 22 0 0 4
658 467
735 467
735 473
766 473
0 1 25 0 0 8192 0 0 22 52 0 3
733 430
733 455
766 455
3 2 25 0 0 4224 0 15 21 0 0 4
660 421
729 421
729 430
763 430
0 6 12 0 0 0 0 0 25 54 0 3
846 190
853 190
853 165
1 5 12 0 0 0 0 25 25 0 0 4
823 165
823 190
847 190
847 165
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
