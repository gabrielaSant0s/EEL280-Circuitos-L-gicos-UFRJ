CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 81 384 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3320 0 0
2
43739.1 10
0
13 Logic Switch~
5 127 385 0 1 11
0 6
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
523 0 0
2
43739.1 9
0
13 Logic Switch~
5 180 385 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 Z1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3557 0 0
2
43739.1 8
0
13 Logic Switch~
5 181 139 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 X1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7246 0 0
2
43739.1 0
0
13 Logic Switch~
5 128 139 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3916 0 0
2
43739.1 0
0
13 Logic Switch~
5 82 138 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
614 0 0
2
43739.1 0
0
9 Inverter~
13 213 178 0 2 22
0 14 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
8494 0 0
2
43739.1 0
0
9 Inverter~
13 215 504 0 2 22
0 7 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
774 0 0
2
43739.1 0
0
9 Inverter~
13 210 442 0 2 22
0 6 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
715 0 0
2
43739.1 0
0
10 2-In NAND~
219 272 433 0 3 22
0 7 4 11
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3281 0 0
2
43739.1 7
0
10 2-In NAND~
219 275 513 0 3 22
0 3 6 9
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3593 0 0
2
43739.1 6
0
10 2-In NAND~
219 411 461 0 3 22
0 11 5 10
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7233 0 0
2
43739.1 3
0
10 2-In NAND~
219 516 486 0 3 22
0 10 9 8
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3410 0 0
2
43739.1 1
0
14 Logic Display~
6 618 466 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3616 0 0
2
43739.1 0
0
14 Logic Display~
6 619 220 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5202 0 0
2
43739.1 0
0
10 2-In NAND~
219 527 241 0 3 22
0 17 16 15
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9145 0 0
2
43739.1 0
0
10 2-In NAND~
219 431 216 0 3 22
0 18 12 17
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9815 0 0
2
43739.1 0
0
9 Inverter~
13 217 276 0 2 22
0 13 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
4766 0 0
2
43739.1 0
0
10 2-In NAND~
219 276 267 0 3 22
0 14 19 16
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8325 0 0
2
43739.1 0
0
10 2-In NAND~
219 273 187 0 3 22
0 2 13 18
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7196 0 0
2
43739.1 0
0
28
2 1 2 0 0 4224 0 7 20 0 0 2
234 178
249 178
2 1 3 0 0 4224 0 8 11 0 0 2
236 504
251 504
2 2 4 0 0 4224 0 9 10 0 0 2
231 442
248 442
1 0 5 0 0 4224 0 3 0 0 0 2
180 397
180 564
1 0 6 0 0 4224 0 2 0 0 0 2
127 397
127 565
1 0 7 0 0 4224 0 1 0 0 0 2
81 396
81 566
3 1 8 0 0 4224 0 13 14 0 0 3
543 486
618 486
618 484
3 2 9 0 0 4224 0 11 13 0 0 4
302 513
464 513
464 495
492 495
3 1 10 0 0 8320 0 12 13 0 0 3
438 461
438 477
492 477
0 2 5 0 0 12416 0 0 12 4 0 4
180 471
195 471
195 470
387 470
3 1 11 0 0 12416 0 10 12 0 0 4
299 433
311 433
311 452
387 452
0 2 6 0 0 0 0 0 11 5 0 2
127 522
251 522
0 1 7 0 0 0 0 0 8 6 0 2
81 504
200 504
0 1 6 0 0 0 0 0 9 5 0 2
127 442
195 442
0 1 7 0 0 0 0 0 10 6 0 2
81 424
248 424
1 0 12 0 0 4224 0 4 0 0 0 2
181 151
181 318
1 0 13 0 0 4224 0 5 0 0 0 2
128 151
128 319
1 0 14 0 0 4224 0 6 0 0 0 2
82 150
82 320
3 1 15 0 0 4224 0 16 15 0 0 3
554 241
619 241
619 238
3 2 16 0 0 4224 0 19 16 0 0 4
303 267
465 267
465 250
503 250
3 1 17 0 0 8320 0 17 16 0 0 3
458 216
458 232
503 232
0 2 12 0 0 4224 0 0 17 16 0 2
181 225
407 225
3 1 18 0 0 12416 0 20 17 0 0 4
300 187
312 187
312 207
407 207
2 2 19 0 0 4224 0 18 19 0 0 2
238 276
252 276
0 1 13 0 0 0 0 0 18 17 0 2
128 276
202 276
1 0 14 0 0 0 0 19 0 0 18 2
252 258
82 258
0 1 14 0 0 128 0 0 7 18 0 2
82 178
198 178
2 0 13 0 0 0 0 20 0 0 17 2
249 196
128 196
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
734 189 971 213
744 197 960 213
27 X = ((X1.(A'B)')' .(AB')')'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
732 450 969 474
742 458 958 474
27 Z = ((Z1.(AB')')' .(A'B)')'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
565 213 590 237
573 221 581 237
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
565 452 590 476
573 460 581 476
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
268 38 481 62
278 46 470 62
24 1)Questao 2 - Comparador
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
