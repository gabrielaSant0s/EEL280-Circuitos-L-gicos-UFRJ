CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 90 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 489
9437202 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 132 130 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3877 0 0
2
43730.1 0
0
13 Logic Switch~
5 182 132 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
926 0 0
2
43730.1 0
0
13 Logic Switch~
5 242 129 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 W
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7262 0 0
2
43730.1 0
0
13 Logic Switch~
5 304 129 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 Z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5267 0 0
2
43730.1 3
0
9 3-In AND~
219 463 523 0 4 22
0 12 11 10 5
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 4 0
1 U
8838 0 0
2
43730.1 0
0
7 Ground~
168 533 434 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7159 0 0
2
43730.1 1
0
4 LED~
171 533 394 0 2 2
10 6 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
5812 0 0
2
43730.1 0
0
9 2-In AND~
219 370 369 0 3 22
0 4 3 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
331 0 0
2
43730.1 2
0
8 2-In OR~
219 438 385 0 3 22
0 9 8 6
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9604 0 0
2
43730.1 1
0
9 2-In AND~
219 369 411 0 3 22
0 7 3 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7518 0 0
2
43730.1 0
0
4 LED~
171 550 532 0 2 2
10 5 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4832 0 0
2
43730.1 1
0
7 Ground~
168 550 572 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6798 0 0
2
43730.1 0
0
8 2-In OR~
219 367 571 0 3 22
0 4 3 10
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3336 0 0
2
43730.1 3
0
8 2-In OR~
219 365 523 0 3 22
0 13 4 11
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8370 0 0
2
43730.1 2
0
8 2-In OR~
219 364 475 0 3 22
0 7 14 12
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3910 0 0
2
43730.1 1
0
7 Ground~
168 597 706 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
316 0 0
2
43730.1 1
0
4 LED~
171 597 662 0 2 2
10 15 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
536 0 0
2
43730.1 0
0
4 LED~
171 543 317 0 2 2
10 16 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4460 0 0
2
43730.1 1
0
7 Ground~
168 543 354 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3260 0 0
2
43730.1 0
0
7 Ground~
168 585 286 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5156 0 0
2
43730.1 0
0
4 LED~
171 585 242 0 2 2
10 17 2
0
0 0 864 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3133 0 0
2
43730.1 0
0
9 3-In AND~
219 371 307 0 4 22
0 13 14 18 16
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
5523 0 0
2
43730.1 0
0
9 2-In AND~
219 372 257 0 3 22
0 7 14 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3746 0 0
2
43730.1 0
0
8 2-In OR~
219 441 231 0 3 22
0 20 19 17
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5668 0 0
2
43730.1 0
0
9 Inverter~
13 99 180 0 2 22
0 14 4
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
5368 0 0
2
43730.1 1
0
9 Inverter~
13 149 182 0 2 22
0 3 18
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
8293 0 0
2
43730.1 1
0
9 Inverter~
13 209 179 0 2 22
0 7 13
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3232 0 0
2
43730.1 1
0
9 Inverter~
13 271 179 0 2 22
0 15 21
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6644 0 0
2
43730.1 2
0
9 2-In AND~
219 373 215 0 3 22
0 14 3 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4978 0 0
2
43730.1 1
0
49
2 0 3 0 0 4096 0 13 0 0 43 2
354 580
182 580
1 0 4 0 0 4096 0 13 0 0 38 2
354 562
102 562
4 1 5 0 0 8320 0 5 11 0 0 3
484 523
484 522
550 522
3 0 6 0 0 4096 0 9 0 0 5 2
471 385
469 385
3 1 6 0 0 12432 0 0 7 0 0 4
465 385
469 385
469 384
533 384
2 1 2 0 0 4112 0 7 6 0 0 2
533 404
533 428
2 0 3 0 0 0 0 10 0 0 43 2
345 420
182 420
1 0 7 0 0 4096 0 10 0 0 46 2
345 402
242 402
2 0 3 0 0 0 0 8 0 0 43 2
346 378
182 378
1 0 4 0 0 0 0 8 0 0 38 2
346 360
102 360
3 2 8 0 0 4224 0 10 9 0 0 4
390 411
417 411
417 394
425 394
3 1 9 0 0 8320 0 8 9 0 0 3
391 369
391 376
425 376
2 1 2 0 0 0 0 11 12 0 0 2
550 542
550 566
3 3 10 0 0 8320 0 13 5 0 0 4
400 571
416 571
416 532
439 532
3 2 11 0 0 4224 0 14 5 0 0 2
398 523
439 523
3 1 12 0 0 8320 0 15 5 0 0 4
397 475
414 475
414 514
439 514
2 0 4 0 0 0 0 14 0 0 38 2
352 532
102 532
1 0 13 0 0 4096 0 14 0 0 44 2
352 514
212 514
2 0 14 0 0 4096 0 15 0 0 40 2
351 484
132 484
1 0 7 0 0 4096 0 15 0 0 46 2
351 466
242 466
3 1 15 0 0 4096 0 0 17 23 0 2
486 652
597 652
2 1 2 0 0 4224 0 17 16 0 0 2
597 672
597 700
0 0 15 0 0 4096 0 0 0 49 21 2
304 652
489 652
4 0 16 0 0 0 0 22 0 0 25 2
392 307
392 307
3 1 16 0 0 8320 0 0 18 0 0 3
388 306
388 307
543 307
2 1 2 0 0 0 0 18 19 0 0 2
543 327
543 348
3 1 17 0 0 8320 0 24 21 0 0 3
474 231
474 232
585 232
2 1 2 0 0 0 0 21 20 0 0 2
585 252
585 280
3 0 18 0 0 4096 0 22 0 0 41 2
347 316
152 316
2 0 14 0 0 0 0 22 0 0 40 2
347 307
132 307
1 0 13 0 0 0 0 22 0 0 44 2
347 298
212 298
3 2 19 0 0 4224 0 23 24 0 0 4
393 257
420 257
420 240
428 240
3 1 20 0 0 8320 0 29 24 0 0 3
394 215
394 222
428 222
2 0 14 0 0 0 0 23 0 0 40 2
348 266
132 266
1 0 7 0 0 0 0 23 0 0 46 2
348 248
242 248
2 0 3 0 0 0 0 29 0 0 43 2
349 224
182 224
1 0 14 0 0 0 0 29 0 0 40 2
349 206
132 206
2 0 4 0 0 4224 0 25 0 0 0 2
102 198
102 756
0 1 14 0 0 0 0 0 25 40 0 3
132 150
102 150
102 162
1 0 14 0 0 4224 0 1 0 0 0 2
132 142
132 757
2 0 18 0 0 4224 0 26 0 0 0 2
152 200
152 758
0 1 3 0 0 0 0 0 26 43 0 3
182 152
152 152
152 164
1 0 3 0 0 4224 0 2 0 0 0 2
182 144
182 759
2 0 13 0 0 4224 0 27 0 0 0 2
212 197
212 755
0 1 7 0 0 0 0 0 27 46 0 3
242 149
212 149
212 161
1 0 7 0 0 4224 0 3 0 0 0 2
242 141
242 756
2 0 21 0 0 4224 0 28 0 0 0 2
274 197
274 755
0 1 15 0 0 0 0 0 28 49 0 3
304 149
274 149
274 161
1 0 15 0 0 4224 0 4 0 0 0 2
304 141
304 756
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
501 492 526 516
509 500 517 516
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
486 609 511 633
494 617 502 633
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
469 355 494 379
477 363 485 379
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
388 277 413 301
396 285 404 301
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
472 186 501 210
482 194 490 210
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
366 18 571 42
376 26 560 42
23 Conversor HEXA para BCD
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
