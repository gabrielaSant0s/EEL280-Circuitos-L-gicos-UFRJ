CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 309 94 0 1 11
0 16
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6187 0 0
2
43737.7 0
0
13 Logic Switch~
5 254 93 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7107 0 0
2
43737.7 0
0
13 Logic Switch~
5 193 93 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6433 0 0
2
43737.7 0
0
13 Logic Switch~
5 126 96 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -30 4 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8559 0 0
2
43737.7 0
0
14 Logic Display~
6 603 477 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3674 0 0
2
43738.7 0
0
10 3-In NAND~
219 527 288 0 4 22
0 5 4 3 20
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
5697 0 0
2
43738.7 0
0
8 2-In OR~
219 495 507 0 3 22
0 7 6 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3805 0 0
2
43738.7 0
0
6 74136~
219 421 575 0 3 22
0 9 8 6
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
5219 0 0
2
43738.7 0
0
6 74136~
219 415 463 0 3 22
0 11 10 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3795 0 0
2
43738.7 0
0
5 4081~
219 358 610 0 3 22
0 13 12 8
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
3637 0 0
2
43738.7 0
0
5 4081~
219 357 549 0 3 22
0 15 14 9
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
3226 0 0
2
43738.7 0
0
5 4081~
219 356 497 0 3 22
0 17 16 10
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
6966 0 0
2
43738.7 0
0
5 4081~
219 355 439 0 3 22
0 19 18 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
9796 0 0
2
43738.7 0
0
14 Logic Display~
6 609 257 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5952 0 0
2
43737.7 0
0
5 7403~
219 420 362 0 3 22
0 21 13 3
0
0 0 624 0
6 74LS38
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3649 0 0
2
43737.7 0
0
5 7403~
219 418 288 0 3 22
0 22 19 4
0
0 0 624 0
6 74LS38
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3716 0 0
2
43737.7 0
0
5 7403~
219 425 203 0 3 22
0 23 18 5
0
0 0 624 0
6 74LS38
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
4797 0 0
2
43737.7 0
0
5 7403~
219 356 353 0 3 22
0 15 16 21
0
0 0 624 0
6 74LS38
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4681 0 0
2
43737.7 0
0
5 7403~
219 354 279 0 3 22
0 14 16 22
0
0 0 624 0
6 74LS38
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9730 0 0
2
43737.7 0
0
5 7403~
219 354 194 0 3 22
0 17 16 23
0
0 0 624 0
6 74LS38
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9874 0 0
2
43737.7 0
0
9 Inverter~
13 292 145 0 2 22
0 16 12
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
364 0 0
2
43737.7 0
0
9 Inverter~
13 236 146 0 2 22
0 17 13
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3656 0 0
2
43737.7 0
0
9 Inverter~
13 174 143 0 2 22
0 14 18
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3131 0 0
2
43737.7 0
0
9 Inverter~
13 106 144 0 2 22
0 15 19
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6772 0 0
2
43737.7 0
0
43
3 1 2 0 0 4224 0 7 5 0 0 3
528 507
603 507
603 495
3 3 3 0 0 8320 0 15 6 0 0 4
447 362
488 362
488 297
503 297
3 2 4 0 0 4224 0 16 6 0 0 2
445 288
503 288
3 1 5 0 0 8320 0 17 6 0 0 4
452 203
493 203
493 279
503 279
3 2 6 0 0 8320 0 8 7 0 0 4
454 575
474 575
474 516
482 516
3 1 7 0 0 8320 0 9 7 0 0 4
448 463
474 463
474 498
482 498
3 2 8 0 0 8320 0 10 8 0 0 4
379 610
397 610
397 584
405 584
3 1 9 0 0 4224 0 11 8 0 0 4
378 549
397 549
397 566
405 566
3 2 10 0 0 8320 0 12 9 0 0 4
377 497
391 497
391 472
399 472
3 1 11 0 0 4224 0 13 9 0 0 4
376 439
391 439
391 454
399 454
2 0 12 0 0 4096 0 10 0 0 35 2
334 619
295 619
1 0 13 0 0 4096 0 10 0 0 34 2
334 601
239 601
2 0 14 0 0 4096 0 11 0 0 42 2
333 558
193 558
1 0 15 0 0 4096 0 11 0 0 43 2
333 540
126 540
2 0 16 0 0 4096 0 12 0 0 40 2
332 506
309 506
1 0 17 0 0 4096 0 12 0 0 41 2
332 488
254 488
2 0 18 0 0 4096 0 13 0 0 33 2
331 448
177 448
1 0 19 0 0 4096 0 13 0 0 32 2
331 430
109 430
4 1 20 0 0 4224 0 6 14 0 0 3
554 288
609 288
609 275
2 0 13 0 0 4096 0 15 0 0 34 2
396 371
239 371
1 3 21 0 0 4224 0 15 18 0 0 2
396 353
383 353
2 0 16 0 0 0 0 18 0 0 40 2
332 362
309 362
1 0 15 0 0 0 0 18 0 0 43 2
332 344
126 344
2 0 19 0 0 4096 0 16 0 0 32 2
394 297
109 297
3 1 22 0 0 4224 0 19 16 0 0 2
381 279
394 279
2 0 16 0 0 0 0 19 0 0 40 2
330 288
309 288
1 0 14 0 0 0 0 19 0 0 42 2
330 270
193 270
2 0 18 0 0 4096 0 17 0 0 33 2
401 212
177 212
3 1 23 0 0 4224 0 20 17 0 0 2
381 194
401 194
2 0 16 0 0 0 0 20 0 0 40 2
330 203
309 203
1 0 17 0 0 0 0 20 0 0 41 2
330 185
254 185
2 0 19 0 0 4224 0 24 0 0 0 2
109 162
109 785
2 0 18 0 0 4224 0 23 0 0 0 2
177 161
177 786
2 0 13 0 0 4224 0 22 0 0 0 2
239 164
239 786
2 0 12 0 0 4224 0 21 0 0 0 2
295 163
295 784
1 0 16 0 0 0 0 21 0 0 40 2
295 127
309 127
1 0 17 0 0 0 0 22 0 0 41 2
239 128
254 128
1 0 14 0 0 0 0 23 0 0 42 2
177 125
193 125
1 0 15 0 0 0 0 24 0 0 43 2
109 126
126 126
1 0 16 0 0 4224 0 1 0 0 0 2
309 106
309 784
1 0 17 0 0 4224 0 2 0 0 0 2
254 105
254 785
1 0 14 0 0 4224 0 3 0 0 0 2
193 105
193 786
1 0 15 0 0 4224 0 4 0 0 0 2
126 108
126 785
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
548 260 577 284
558 268 566 284
1 M
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
