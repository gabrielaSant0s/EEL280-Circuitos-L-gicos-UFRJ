CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 140 240 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 140 170 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89908e-315 0
0
5 4011~
219 312 231 0 3 22
0 6 7 4
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 3 0
1 U
3124 0 0
2
5.89908e-315 0
0
5 4011~
219 402 200 0 3 22
0 5 4 3
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 3 0
1 U
3421 0 0
2
5.89908e-315 0
0
5 4011~
219 311 179 0 3 22
0 8 6 5
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 3 0
1 U
8157 0 0
2
5.89908e-315 0
0
5 4011~
219 222 203 0 3 22
0 8 7 6
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
5.89908e-315 0
0
7 Ground~
168 481 267 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
5.89908e-315 0
0
4 LED~
171 481 227 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7361 0 0
2
5.89908e-315 0
0
10
2 1 2 0 0 4224 0 8 7 0 0 2
481 237
481 261
3 1 3 0 0 4224 0 4 8 0 0 3
429 200
481 200
481 217
3 2 4 0 0 8320 0 3 4 0 0 4
339 231
358 231
358 209
378 209
3 1 5 0 0 4224 0 5 4 0 0 4
338 179
358 179
358 191
378 191
0 1 6 0 0 8320 0 0 3 6 0 3
268 203
268 222
288 222
3 2 6 0 0 0 0 6 5 0 0 4
249 203
269 203
269 188
287 188
0 2 7 0 0 4224 0 0 3 9 0 2
191 240
288 240
0 1 8 0 0 4224 0 0 5 10 0 2
191 170
287 170
1 2 7 0 0 0 0 1 6 0 0 4
152 240
191 240
191 212
198 212
1 1 8 0 0 0 0 2 6 0 0 4
152 170
191 170
191 194
198 194
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 114
610 122 895 226
620 130 884 210
114 A B | A xor B | ( A'+B' ).( A+B ) 
0 0 |   0     |		0
0 1 |   1     |		1
1 0 |   1     |		1
1 1 |   0     |		0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
