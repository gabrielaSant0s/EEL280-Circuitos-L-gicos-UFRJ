CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1380 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.168350
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
111
13 Logic Switch~
5 950 2726 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 x1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9597 0 0
2
43729.2 3
0
13 Logic Switch~
5 1006 2726 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 y1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9950 0 0
2
43729.2 2
0
13 Logic Switch~
5 1056 2725 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 w1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3239 0 0
2
43729.2 1
0
13 Logic Switch~
5 1107 2723 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 z1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7621 0 0
2
43729.2 0
0
13 Logic Switch~
5 246 1459 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8673 0 0
2
5.89909e-315 5.38788e-315
0
13 Logic Switch~
5 195 1461 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 w
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9712 0 0
2
5.89909e-315 5.39306e-315
0
13 Logic Switch~
5 145 1462 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3900 0 0
2
5.89909e-315 5.39824e-315
0
13 Logic Switch~
5 89 1462 0 1 11
0 28
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 x
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4153 0 0
2
5.89909e-315 5.40342e-315
0
13 Logic Switch~
5 290 85 0 1 11
0 94
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8251 0 0
2
43729.1 0
0
13 Logic Switch~
5 226 83 0 1 11
0 77
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 W
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8341 0 0
2
43729.1 1
0
13 Logic Switch~
5 174 82 0 1 11
0 79
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6192 0 0
2
43729.1 2
0
13 Logic Switch~
5 116 82 0 1 11
0 82
0
0 0 21360 270
2 0V
-7 -21 7 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3842 0 0
2
43729.1 3
0
9 Inverter~
13 985 2784 0 2 22
0 8 105
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U34E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 5 36 0
1 U
6185 0 0
2
43729.2 7
0
9 Inverter~
13 920 2783 0 2 22
0 9 106
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U34D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 4 36 0
1 U
3914 0 0
2
43729.2 6
0
9 Inverter~
13 1086 2790 0 2 22
0 6 107
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U34C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 3 36 0
1 U
367 0 0
2
43729.2 5
0
9 Inverter~
13 1036 2789 0 2 22
0 7 108
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U34B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 2 36 0
1 U
4366 0 0
2
43729.2 4
0
9 2-In AND~
219 358 2827 0 3 22
0 10 4 32
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U40D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 42 0
1 U
7433 0 0
2
43729.2 0
0
7 Ground~
168 950 2040 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8588 0 0
2
43729.2 0
0
9 CC 7-Seg~
183 864 1875 0 17 19
10 12 18 17 16 15 14 13 109 2
1 0 1 1 1 1 1 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6897 0 0
2
43729.2 0
0
9 2-In AND~
219 320 2920 0 3 22
0 28 26 23
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U36D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 38 0
1 U
3458 0 0
2
43729.2 7
0
9 2-In AND~
219 319 2973 0 3 22
0 27 10 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U40A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 42 0
1 U
5508 0 0
2
43729.2 6
0
9 2-In AND~
219 319 3018 0 3 22
0 11 28 25
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U40B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 42 0
1 U
3981 0 0
2
43729.2 5
0
9 2-In AND~
219 320 3065 0 3 22
0 27 26 24
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U40C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 42 0
1 U
4581 0 0
2
43729.2 4
0
9 3-In AND~
219 321 3107 0 4 22
0 3 5 4 19
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U37B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 39 0
1 U
3346 0 0
2
43729.2 3
0
8 2-In OR~
219 402 2937 0 3 22
0 23 22 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U39B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 41 0
1 U
8843 0 0
2
43729.2 2
0
8 2-In OR~
219 401 3038 0 3 22
0 25 24 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U39C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 41 0
1 U
566 0 0
2
43729.2 1
0
8 3-In OR~
219 502 3038 0 4 22
0 21 20 19 13
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U38B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 40 0
1 U
3750 0 0
2
43729.2 0
0
9 2-In AND~
219 359 2700 0 3 22
0 3 10 35
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U36A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 38 0
1 U
9887 0 0
2
43729.1 7
0
9 2-In AND~
219 359 2742 0 3 22
0 28 26 34
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U36B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 38 0
1 U
351 0 0
2
43729.1 6
0
9 2-In AND~
219 359 2784 0 3 22
0 27 28 33
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U36C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 38 0
1 U
7542 0 0
2
43729.1 5
0
9 3-In AND~
219 357 2869 0 4 22
0 5 4 3 31
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U37A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 39 0
1 U
9283 0 0
2
43729.1 3
0
8 3-In OR~
219 438 2720 0 4 22
0 35 34 33 30
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U38A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 40 0
1 U
3600 0 0
2
43729.1 2
0
8 2-In OR~
219 445 2819 0 3 22
0 32 31 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 21 0
1 U
8274 0 0
2
43729.1 1
0
8 2-In OR~
219 530 2764 0 3 22
0 30 29 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U39A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 41 0
1 U
3329 0 0
2
43729.1 0
0
9 2-In AND~
219 367 2548 0 3 22
0 28 4 40
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 35 0
1 U
3509 0 0
2
43729.1 5
0
9 4-In NOR~
219 464 2597 0 5 22
0 40 39 38 37 36
0
0 0 624 0
4 4002
-14 -24 14 -16
4 U35A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 37 0
1 U
90 0 0
2
43729.1 4
0
9 2-In AND~
219 369 2585 0 3 22
0 27 10 39
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 35 0
1 U
5259 0 0
2
43729.1 3
0
9 2-In AND~
219 369 2624 0 3 22
0 26 10 38
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 35 0
1 U
6548 0 0
2
43729.1 2
0
9 2-In AND~
219 369 2663 0 3 22
0 28 27 37
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U33D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 35 0
1 U
9326 0 0
2
43729.1 1
0
9 Inverter~
13 541 2597 0 2 22
0 36 15
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U34A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 36 0
1 U
5634 0 0
2
43729.1 0
0
9 2-In AND~
219 417 2333 0 3 22
0 3 28 47
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U28D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
7902 0 0
2
5.89909e-315 5.37752e-315
0
9 3-In AND~
219 418 2426 0 4 22
0 10 5 26 45
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U26B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 28 0
1 U
6805 0 0
2
5.89909e-315 5.36716e-315
0
9 3-In AND~
219 419 2470 0 4 22
0 27 11 26 43
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U26C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 28 0
1 U
6198 0 0
2
5.89909e-315 5.3568e-315
0
9 3-In AND~
219 420 2514 0 4 22
0 3 11 4 44
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U32A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 34 0
1 U
9216 0 0
2
5.89909e-315 5.34643e-315
0
9 3-In AND~
219 417 2382 0 4 22
0 27 10 4 46
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U32B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 34 0
1 U
9719 0 0
2
5.89909e-315 5.32571e-315
0
8 2-In OR~
219 485 2348 0 3 22
0 47 46 42
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
3781 0 0
2
5.89909e-315 5.30499e-315
0
8 2-In OR~
219 578 2411 0 3 22
0 42 41 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 21 0
1 U
8277 0 0
2
5.89909e-315 5.26354e-315
0
8 3-In OR~
219 501 2469 0 4 22
0 45 43 44 41
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 10 0
1 U
3457 0 0
2
5.89909e-315 0
0
9 2-In XOR~
219 301 2143 0 3 22
0 28 4 51
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U29B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
3796 0 0
2
5.89909e-315 5.3568e-315
0
9 2-In AND~
219 309 2208 0 3 22
0 3 11 50
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U28B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
6904 0 0
2
5.89909e-315 5.34643e-315
0
10 2-In NAND~
219 311 2276 0 3 22
0 27 10 52
0
0 0 624 0
6 74LS37
-14 -24 28 -16
4 U27C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 29 0
1 U
8602 0 0
2
5.89909e-315 5.32571e-315
0
9 2-In AND~
219 385 2294 0 3 22
0 52 5 48
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U28C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
3607 0 0
2
5.89909e-315 5.30499e-315
0
8 2-In OR~
219 393 2170 0 3 22
0 51 50 49
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U25D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
9456 0 0
2
5.89909e-315 5.26354e-315
0
8 2-In OR~
219 485 2233 0 3 22
0 49 48 17
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U30A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
3348 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 560 2025 0 3 22
0 53 54 18
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U25C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
7418 0 0
2
5.89909e-315 5.36716e-315
0
8 2-In OR~
219 466 1932 0 3 22
0 56 55 53
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U25B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 27 0
1 U
3281 0 0
2
5.89909e-315 5.3568e-315
0
9 2-In AND~
219 379 2103 0 3 22
0 57 26 54
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U28A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
3613 0 0
2
5.89909e-315 5.34643e-315
0
10 2-In NAND~
219 312 2060 0 3 22
0 28 11 57
0
0 0 624 0
6 74LS37
-14 -24 28 -16
4 U27A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
9506 0 0
2
5.89909e-315 5.32571e-315
0
9 2-In AND~
219 392 1986 0 3 22
0 58 5 55
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U21D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 23 0
1 U
6773 0 0
2
5.89909e-315 5.30499e-315
0
6 74266~
219 302 1949 0 3 22
0 27 11 58
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
8799 0 0
2
5.89909e-315 5.26354e-315
0
9 3-In AND~
219 320 1886 0 4 22
0 28 3 11 56
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U26A
-20 18 8 26
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 28 0
1 U
7433 0 0
2
5.89909e-315 0
0
7 Ground~
168 1422 1643 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6183 0 0
2
5.89909e-315 5.26354e-315
0
4 LED~
171 1422 1611 0 2 2
10 59 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5243 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 610 1711 0 3 22
0 60 61 12
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U22D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 24 0
1 U
3217 0 0
2
5.89909e-315 5.44487e-315
0
8 2-In OR~
219 520 1632 0 3 22
0 63 62 60
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U22B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 24 0
1 U
998 0 0
2
5.89909e-315 5.44746e-315
0
8 2-In OR~
219 444 1821 0 3 22
0 65 64 61
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U22A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
9272 0 0
2
5.89909e-315 5.45005e-315
0
8 2-In OR~
219 436 1701 0 3 22
0 67 66 62
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
3327 0 0
2
5.89909e-315 5.45264e-315
0
8 2-In OR~
219 427 1583 0 3 22
0 69 68 63
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
466 0 0
2
5.89909e-315 5.45523e-315
0
9 3-In AND~
219 320 1847 0 4 22
0 28 26 3 64
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 18 0
1 U
6854 0 0
2
5.89909e-315 5.45782e-315
0
9 3-In AND~
219 321 1793 0 4 22
0 11 5 4 65
0
0 0 624 0
5 74F11
-18 -28 17 -20
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 18 0
1 U
7745 0 0
2
5.89909e-315 5.46041e-315
0
9 2-In AND~
219 324 1729 0 3 22
0 10 26 66
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 23 0
1 U
5764 0 0
2
5.89909e-315 5.463e-315
0
9 2-In AND~
219 324 1671 0 3 22
0 28 10 67
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5379 0 0
2
5.89909e-315 5.46559e-315
0
9 2-In AND~
219 324 1615 0 3 22
0 4 27 68
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7186 0 0
2
5.89909e-315 5.46818e-315
0
9 2-In AND~
219 322 1553 0 3 22
0 5 27 69
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9136 0 0
2
5.89909e-315 5.47077e-315
0
9 Inverter~
13 175 1525 0 2 22
0 27 3
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U20A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 22 0
1 U
7143 0 0
2
5.89909e-315 5.47207e-315
0
9 Inverter~
13 225 1526 0 2 22
0 11 10
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
9634 0 0
2
5.89909e-315 5.47336e-315
0
9 Inverter~
13 59 1519 0 2 22
0 28 5
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
3661 0 0
2
5.89909e-315 5.47466e-315
0
9 Inverter~
13 124 1520 0 2 22
0 4 26
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U10D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
4323 0 0
2
5.89909e-315 5.47595e-315
0
7 Ground~
168 674 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9804 0 0
2
5.89909e-315 5.48502e-315
0
9 CC 7-Seg~
183 607 384 0 17 19
10 76 75 74 73 72 71 70 110 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3981 0 0
2
5.89909e-315 5.48631e-315
0
8 2-In OR~
219 515 1013 0 3 22
0 82 84 87
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
9102 0 0
2
5.89909e-315 5.48761e-315
0
8 2-In OR~
219 508 1124 0 3 22
0 86 85 83
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
6812 0 0
2
5.89909e-315 5.4889e-315
0
8 2-In OR~
219 579 1073 0 3 22
0 87 83 70
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
6462 0 0
2
5.89909e-315 5.4902e-315
0
9 2-In AND~
219 416 1034 0 3 22
0 77 78 84
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
5184 0 0
2
5.89909e-315 5.49149e-315
0
9 2-In AND~
219 416 1092 0 3 22
0 79 80 86
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
9835 0 0
2
5.89909e-315 5.49279e-315
0
9 2-In AND~
219 415 1151 0 3 22
0 77 81 85
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
8927 0 0
2
5.89909e-315 5.49408e-315
0
8 2-In OR~
219 557 892 0 3 22
0 89 88 71
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3701 0 0
2
5.89909e-315 5.49538e-315
0
8 2-In OR~
219 482 930 0 3 22
0 91 90 88
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
5444 0 0
2
5.89909e-315 5.49667e-315
0
8 2-In OR~
219 485 855 0 3 22
0 92 82 89
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
4858 0 0
2
5.89909e-315 5.49797e-315
0
9 2-In AND~
219 409 832 0 3 22
0 79 81 92
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
4290 0 0
2
5.89909e-315 5.49926e-315
0
9 2-In AND~
219 408 899 0 3 22
0 79 80 91
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
4394 0 0
2
5.89909e-315 5.50056e-315
0
9 2-In AND~
219 405 958 0 3 22
0 80 81 90
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
7544 0 0
2
5.89909e-315 5.50185e-315
0
9 2-In AND~
219 553 746 0 3 22
0 93 81 72
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
5696 0 0
2
5.89909e-315 5.50315e-315
0
8 2-In OR~
219 446 717 0 3 22
0 78 77 93
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
5601 0 0
2
5.89909e-315 5.50444e-315
0
9 3-In AND~
219 399 636 0 4 22
0 80 94 79 97
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 6 0
1 U
4406 0 0
2
43729.1 4
0
8 3-In OR~
219 556 553 0 4 22
0 99 98 97 73
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
882 0 0
2
43729.1 5
0
8 3-In OR~
219 485 470 0 4 22
0 82 96 95 99
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
3359 0 0
2
43729.1 6
0
9 2-In AND~
219 403 481 0 3 22
0 81 77 96
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4933 0 0
2
43729.1 7
0
9 2-In AND~
219 402 530 0 3 22
0 78 81 95
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
9209 0 0
2
43729.1 8
0
9 2-In AND~
219 397 588 0 3 22
0 78 77 98
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
7797 0 0
2
43729.1 9
0
8 2-In OR~
219 495 385 0 3 22
0 79 100 74
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
6403 0 0
2
43729.1 10
0
8 2-In OR~
219 412 411 0 3 22
0 80 94 100
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3709 0 0
2
43729.1 11
0
6 74266~
219 369 352 0 3 22
0 77 94 101
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9784 0 0
2
43729.1 12
0
8 2-In OR~
219 491 303 0 3 22
0 78 101 75
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6816 0 0
2
43729.1 13
0
8 2-In OR~
219 388 188 0 3 22
0 82 77 103
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7493 0 0
2
43729.1 14
0
8 2-In OR~
219 485 221 0 3 22
0 103 102 76
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5587 0 0
2
43729.1 15
0
6 74266~
219 390 264 0 3 22
0 79 94 102
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
5642 0 0
2
43729.1 16
0
9 Inverter~
13 260 136 0 2 22
0 94 81
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
3577 0 0
2
43729.1 17
0
9 Inverter~
13 199 134 0 2 22
0 77 80
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
3255 0 0
2
43729.1 18
0
9 Inverter~
13 143 131 0 2 22
0 79 78
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
345 0 0
2
43729.1 19
0
9 Inverter~
13 82 132 0 2 22
0 82 104
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3918 0 0
2
43729.1 20
0
230
3 0 3 0 0 4096 0 31 0 0 143 2
333 2878
178 2878
2 0 4 0 0 4096 0 31 0 0 151 2
333 2869
145 2869
1 0 5 0 0 4096 0 31 0 0 141 2
333 2860
62 2860
1 0 6 0 0 4112 0 15 0 0 8 3
1089 2772
1089 2747
1107 2747
1 0 7 0 0 4112 0 16 0 0 9 3
1039 2771
1039 2747
1056 2747
1 0 8 0 0 4112 0 13 0 0 10 3
988 2766
988 2748
1006 2748
1 0 9 0 0 8208 0 14 0 0 11 3
923 2765
923 2750
950 2750
1 0 6 0 0 4240 0 4 0 0 0 2
1107 2735
1107 4529
1 0 7 0 0 4240 0 3 0 0 0 2
1056 2737
1056 4528
1 0 8 0 0 4240 0 2 0 0 0 2
1006 2738
1006 4528
1 0 9 0 0 4240 0 1 0 0 0 2
950 2738
950 4528
2 0 4 0 0 4096 0 17 0 0 151 2
334 2836
145 2836
1 0 10 0 0 4096 0 17 0 0 144 2
334 2818
228 2818
1 0 11 0 0 4096 0 22 0 0 149 2
295 3009
246 3009
9 1 2 0 0 8320 0 19 18 0 0 3
864 1833
950 1833
950 2034
3 1 12 0 0 8320 0 64 19 0 0 5
643 1711
758 1711
758 1921
843 1921
843 1911
7 4 13 0 0 4224 0 19 27 0 0 3
879 1911
879 3038
535 3038
6 3 14 0 0 4224 0 19 34 0 0 3
873 1911
873 2764
563 2764
5 2 15 0 0 4224 0 19 40 0 0 3
867 1911
867 2597
562 2597
4 3 16 0 0 4224 0 19 47 0 0 3
861 1911
861 2411
611 2411
3 3 17 0 0 4224 0 54 19 0 0 3
518 2233
855 2233
855 1911
3 2 18 0 0 12416 0 55 19 0 0 5
593 2025
709 2025
709 2043
849 2043
849 1911
4 3 19 0 0 4224 0 24 27 0 0 4
342 3107
465 3107
465 3047
489 3047
3 2 20 0 0 4224 0 26 27 0 0 2
434 3038
490 3038
3 1 21 0 0 8320 0 25 27 0 0 4
435 2937
464 2937
464 3029
489 3029
3 2 22 0 0 4224 0 21 25 0 0 4
340 2973
367 2973
367 2946
389 2946
3 1 23 0 0 4224 0 20 25 0 0 4
341 2920
367 2920
367 2928
389 2928
3 2 24 0 0 4224 0 23 26 0 0 4
341 3065
369 3065
369 3047
388 3047
3 1 25 0 0 4224 0 22 26 0 0 4
340 3018
368 3018
368 3029
388 3029
3 0 4 0 0 0 0 24 0 0 151 2
297 3116
145 3116
2 0 5 0 0 0 0 24 0 0 141 2
297 3107
62 3107
1 0 3 0 0 0 0 24 0 0 143 2
297 3098
178 3098
2 0 26 0 0 4096 0 23 0 0 142 2
296 3074
127 3074
1 0 27 0 0 4096 0 23 0 0 150 2
296 3056
195 3056
2 0 28 0 0 4096 0 22 0 0 152 2
295 3027
89 3027
2 0 10 0 0 0 0 21 0 0 144 2
295 2982
228 2982
1 0 27 0 0 0 0 21 0 0 150 2
295 2964
195 2964
2 0 26 0 0 0 0 20 0 0 142 2
296 2929
127 2929
1 0 28 0 0 4096 0 20 0 0 152 2
296 2911
89 2911
3 2 29 0 0 8320 0 33 34 0 0 4
478 2819
489 2819
489 2773
517 2773
4 1 30 0 0 8320 0 32 34 0 0 4
471 2720
488 2720
488 2755
517 2755
4 2 31 0 0 8320 0 31 33 0 0 4
378 2869
416 2869
416 2828
432 2828
3 1 32 0 0 8320 0 17 33 0 0 3
379 2827
379 2810
432 2810
3 3 33 0 0 8320 0 30 32 0 0 4
380 2784
416 2784
416 2729
425 2729
3 2 34 0 0 12416 0 29 32 0 0 4
380 2742
398 2742
398 2720
426 2720
3 1 35 0 0 12416 0 28 32 0 0 4
380 2700
399 2700
399 2711
425 2711
2 0 28 0 0 4096 0 30 0 0 152 2
335 2793
89 2793
1 0 27 0 0 4096 0 30 0 0 150 2
335 2775
195 2775
2 0 26 0 0 4096 0 29 0 0 142 2
335 2751
127 2751
1 0 28 0 0 0 0 29 0 0 152 2
335 2733
89 2733
2 0 10 0 0 4096 0 28 0 0 144 2
335 2709
228 2709
1 0 3 0 0 4096 0 28 0 0 143 2
335 2691
178 2691
2 0 10 0 0 4096 0 37 0 0 144 2
345 2594
228 2594
5 0 36 0 0 0 0 36 0 0 55 2
503 2597
503 2597
3 1 36 0 0 4224 0 0 40 0 0 2
498 2597
526 2597
3 4 37 0 0 8320 0 39 36 0 0 4
390 2663
436 2663
436 2611
447 2611
3 3 38 0 0 12416 0 38 36 0 0 4
390 2624
415 2624
415 2602
447 2602
3 2 39 0 0 8320 0 37 36 0 0 3
390 2585
390 2593
447 2593
3 1 40 0 0 8320 0 35 36 0 0 4
388 2548
413 2548
413 2584
447 2584
2 0 27 0 0 4096 0 39 0 0 150 2
345 2672
195 2672
1 0 28 0 0 4096 0 39 0 0 152 2
345 2654
89 2654
2 0 10 0 0 0 0 38 0 0 144 2
345 2633
228 2633
1 0 26 0 0 4096 0 38 0 0 142 2
345 2615
127 2615
1 0 27 0 0 0 0 37 0 0 150 2
345 2576
195 2576
2 0 4 0 0 4096 0 35 0 0 151 2
343 2557
145 2557
1 0 28 0 0 0 0 35 0 0 152 2
343 2539
89 2539
2 0 11 0 0 4096 0 44 0 0 149 2
396 2514
246 2514
4 2 41 0 0 8320 0 48 47 0 0 4
534 2469
538 2469
538 2420
565 2420
3 1 42 0 0 8320 0 46 47 0 0 4
518 2348
538 2348
538 2402
565 2402
4 2 43 0 0 4224 0 43 48 0 0 4
440 2470
482 2470
482 2469
489 2469
4 3 44 0 0 8320 0 44 48 0 0 4
441 2514
472 2514
472 2478
488 2478
4 1 45 0 0 8320 0 42 48 0 0 4
439 2426
455 2426
455 2460
488 2460
4 2 46 0 0 8320 0 45 46 0 0 4
438 2382
455 2382
455 2357
472 2357
3 1 47 0 0 12416 0 41 46 0 0 4
438 2333
451 2333
451 2339
472 2339
3 0 4 0 0 4096 0 44 0 0 151 2
396 2523
145 2523
1 0 3 0 0 4096 0 44 0 0 143 2
396 2505
178 2505
3 0 26 0 0 4096 0 43 0 0 142 2
395 2479
127 2479
2 0 11 0 0 128 0 43 0 0 149 2
395 2470
246 2470
1 0 27 0 0 4096 0 43 0 0 150 2
395 2461
195 2461
3 0 26 0 0 0 0 42 0 0 142 2
394 2435
127 2435
2 0 5 0 0 4096 0 42 0 0 141 2
394 2426
62 2426
1 0 10 0 0 4096 0 42 0 0 144 2
394 2417
228 2417
3 0 4 0 0 0 0 45 0 0 151 2
393 2391
145 2391
2 0 10 0 0 0 0 45 0 0 144 2
393 2382
228 2382
1 0 27 0 0 0 0 45 0 0 150 2
393 2373
195 2373
2 0 28 0 0 4096 0 41 0 0 152 2
393 2342
89 2342
1 0 3 0 0 0 0 41 0 0 143 2
393 2324
178 2324
3 2 48 0 0 4224 0 52 54 0 0 4
406 2294
464 2294
464 2242
472 2242
3 1 49 0 0 8320 0 53 54 0 0 4
426 2170
464 2170
464 2224
472 2224
3 2 50 0 0 4224 0 50 53 0 0 4
330 2208
372 2208
372 2179
380 2179
3 1 51 0 0 4224 0 49 53 0 0 4
334 2143
372 2143
372 2161
380 2161
2 0 5 0 0 0 0 52 0 0 141 2
361 2303
62 2303
3 1 52 0 0 4224 0 51 52 0 0 4
338 2276
353 2276
353 2285
361 2285
1 0 27 0 0 0 0 51 0 0 150 2
287 2267
195 2267
2 0 10 0 0 0 0 51 0 0 144 2
287 2285
228 2285
2 0 11 0 0 0 0 50 0 0 149 2
285 2217
246 2217
1 0 3 0 0 0 0 50 0 0 143 2
285 2199
178 2199
2 0 4 0 0 0 0 49 0 0 151 2
285 2152
145 2152
1 0 28 0 0 0 0 49 0 0 152 2
285 2134
89 2134
3 1 53 0 0 8320 0 56 55 0 0 4
499 1932
526 1932
526 2016
547 2016
3 2 54 0 0 4224 0 57 55 0 0 4
400 2103
526 2103
526 2034
547 2034
3 2 55 0 0 8320 0 59 56 0 0 4
413 1986
439 1986
439 1941
453 1941
4 1 56 0 0 4224 0 61 56 0 0 4
341 1886
439 1886
439 1923
453 1923
2 0 26 0 0 0 0 57 0 0 142 2
355 2112
127 2112
3 1 57 0 0 8320 0 58 57 0 0 4
339 2060
347 2060
347 2094
355 2094
2 0 11 0 0 0 0 58 0 0 149 2
288 2069
246 2069
1 0 28 0 0 0 0 58 0 0 152 2
288 2051
89 2051
2 0 5 0 0 0 0 59 0 0 141 2
368 1995
62 1995
3 1 58 0 0 8320 0 60 59 0 0 4
341 1949
360 1949
360 1977
368 1977
2 0 11 0 0 0 0 60 0 0 149 2
286 1958
246 1958
1 0 27 0 0 0 0 60 0 0 150 2
286 1940
195 1940
3 0 11 0 0 0 0 61 0 0 149 2
296 1895
246 1895
2 0 3 0 0 0 0 61 0 0 143 2
296 1886
178 1886
1 0 28 0 0 0 0 61 0 0 152 2
296 1877
89 1877
3 1 59 0 0 4224 0 0 63 0 0 3
1385 1572
1422 1572
1422 1601
1 2 2 0 0 0 0 62 63 0 0 2
1422 1637
1422 1621
3 1 60 0 0 8320 0 65 64 0 0 4
553 1632
589 1632
589 1702
597 1702
3 2 61 0 0 8320 0 66 64 0 0 4
477 1821
563 1821
563 1720
597 1720
3 2 62 0 0 8320 0 67 65 0 0 4
469 1701
499 1701
499 1641
507 1641
3 1 63 0 0 8320 0 68 65 0 0 4
460 1583
499 1583
499 1623
507 1623
4 2 64 0 0 4224 0 69 66 0 0 4
341 1847
423 1847
423 1830
431 1830
4 1 65 0 0 4224 0 70 66 0 0 4
342 1793
423 1793
423 1812
431 1812
3 2 66 0 0 4224 0 71 67 0 0 4
345 1729
417 1729
417 1710
423 1710
3 1 67 0 0 4224 0 72 67 0 0 4
345 1671
417 1671
417 1692
423 1692
3 2 68 0 0 4224 0 73 68 0 0 4
345 1615
407 1615
407 1592
414 1592
3 1 69 0 0 4224 0 74 68 0 0 4
343 1553
407 1553
407 1574
414 1574
3 0 3 0 0 0 0 69 0 0 143 2
296 1856
178 1856
2 0 26 0 0 0 0 69 0 0 142 2
296 1847
127 1847
1 0 28 0 0 0 0 72 0 0 152 2
300 1662
89 1662
1 0 28 0 0 0 0 69 0 0 152 2
296 1838
89 1838
3 0 4 0 0 0 0 70 0 0 151 2
297 1802
145 1802
2 0 5 0 0 0 0 70 0 0 141 2
297 1793
62 1793
1 0 11 0 0 0 0 70 0 0 149 2
297 1784
246 1784
2 0 26 0 0 0 0 71 0 0 142 2
300 1738
127 1738
1 0 10 0 0 0 0 71 0 0 144 2
300 1720
228 1720
2 0 10 0 0 0 0 72 0 0 144 2
300 1680
228 1680
2 0 27 0 0 0 0 73 0 0 150 2
300 1624
195 1624
1 0 4 0 0 0 0 73 0 0 151 2
300 1606
145 1606
2 0 27 0 0 0 0 74 0 0 150 2
298 1562
195 1562
0 1 5 0 0 0 0 0 74 141 0 3
62 1543
62 1544
298 1544
2 0 5 0 0 4224 0 77 0 0 0 2
62 1537
62 3263
2 0 26 0 0 4224 0 78 0 0 0 2
127 1538
127 3262
2 0 3 0 0 4224 0 75 0 0 0 2
178 1543
178 3263
2 0 10 0 0 4224 0 76 0 0 0 2
228 1544
228 3264
1 0 11 0 0 0 0 76 0 0 149 3
228 1508
228 1483
246 1483
1 0 27 0 0 0 0 75 0 0 150 3
178 1507
178 1483
195 1483
1 0 4 0 0 0 0 78 0 0 151 3
127 1502
127 1484
145 1484
1 0 28 0 0 0 0 77 0 0 152 3
62 1501
62 1486
89 1486
1 0 11 0 0 4224 0 5 0 0 0 2
246 1471
246 3265
1 0 27 0 0 4224 0 6 0 0 0 2
195 1473
195 3264
1 0 4 0 0 4224 0 7 0 0 0 2
145 1474
145 3264
1 0 28 0 0 4224 0 8 0 0 0 2
89 1474
89 3264
7 3 70 0 0 4224 0 80 83 0 0 3
622 420
622 1073
612 1073
6 3 71 0 0 4224 0 80 87 0 0 3
616 420
616 892
590 892
5 3 72 0 0 4224 0 80 93 0 0 3
610 420
610 746
574 746
4 4 73 0 0 4224 0 80 96 0 0 3
604 420
604 553
589 553
3 3 74 0 0 8320 0 80 101 0 0 5
598 420
598 430
541 430
541 385
528 385
2 3 75 0 0 12416 0 80 104 0 0 5
592 420
592 425
537 425
537 303
524 303
1 3 76 0 0 8320 0 80 106 0 0 4
586 420
533 420
533 221
518 221
1 9 2 0 0 128 0 79 80 0 0 4
674 426
674 330
607 330
607 342
1 0 77 0 0 4096 0 84 0 0 223 2
392 1025
226 1025
2 0 78 0 0 4096 0 84 0 0 226 2
392 1043
146 1043
1 0 79 0 0 4096 0 85 0 0 227 2
392 1083
174 1083
2 0 80 0 0 4096 0 85 0 0 222 2
392 1101
202 1101
2 0 81 0 0 4096 0 86 0 0 220 2
391 1160
263 1160
1 0 77 0 0 0 0 86 0 0 223 2
391 1142
226 1142
1 0 82 0 0 4096 0 81 0 0 230 2
502 1004
116 1004
3 2 83 0 0 8320 0 82 83 0 0 4
541 1124
558 1124
558 1082
566 1082
3 2 84 0 0 4224 0 84 81 0 0 4
437 1034
471 1034
471 1022
502 1022
3 2 85 0 0 4224 0 86 82 0 0 4
436 1151
476 1151
476 1133
495 1133
3 1 86 0 0 4224 0 85 82 0 0 4
437 1092
476 1092
476 1115
495 1115
3 1 87 0 0 4224 0 81 83 0 0 3
548 1013
548 1064
566 1064
2 0 81 0 0 0 0 92 0 0 220 2
381 967
263 967
2 0 80 0 0 0 0 91 0 0 222 2
384 908
202 908
1 0 80 0 0 0 0 92 0 0 222 2
381 949
202 949
2 0 81 0 0 0 0 90 0 0 220 2
385 841
263 841
1 0 79 0 0 0 0 90 0 0 227 2
385 823
174 823
2 0 82 0 0 0 0 89 0 0 230 2
472 864
116 864
3 2 88 0 0 8320 0 88 87 0 0 4
515 930
536 930
536 901
544 901
3 1 89 0 0 8320 0 89 87 0 0 4
518 855
536 855
536 883
544 883
3 2 90 0 0 4224 0 92 88 0 0 4
426 958
461 958
461 939
469 939
3 1 91 0 0 4224 0 91 88 0 0 4
429 899
461 899
461 921
469 921
3 1 92 0 0 8320 0 90 89 0 0 3
430 832
430 846
472 846
0 1 79 0 0 0 0 0 91 227 0 2
174 890
384 890
0 2 81 0 0 4096 0 0 93 220 0 4
263 781
513 781
513 755
529 755
3 1 93 0 0 4224 0 94 93 0 0 4
479 717
512 717
512 737
529 737
0 2 77 0 0 4096 0 0 94 223 0 4
226 741
396 741
396 726
433 726
0 1 78 0 0 4096 0 0 94 226 0 4
146 693
396 693
396 708
433 708
3 0 79 0 0 0 0 95 0 0 227 2
375 645
174 645
2 0 94 0 0 4096 0 95 0 0 219 2
375 636
290 636
1 0 80 0 0 0 0 95 0 0 222 2
375 627
202 627
2 0 77 0 0 0 0 100 0 0 223 2
373 597
226 597
1 0 78 0 0 0 0 100 0 0 226 2
373 579
146 579
2 0 81 0 0 0 0 99 0 0 220 2
378 539
263 539
1 0 81 0 0 0 0 98 0 0 220 2
379 472
263 472
1 0 78 0 0 0 0 99 0 0 226 2
378 521
146 521
2 0 77 0 0 0 0 98 0 0 223 2
379 490
226 490
3 3 95 0 0 8320 0 99 97 0 0 4
423 530
452 530
452 479
472 479
3 2 96 0 0 12416 0 98 97 0 0 4
424 481
440 481
440 470
473 470
1 0 82 0 0 0 0 97 0 0 230 2
472 461
116 461
4 3 97 0 0 4224 0 95 96 0 0 4
420 636
520 636
520 562
543 562
3 2 98 0 0 4224 0 100 96 0 0 4
418 588
495 588
495 553
544 553
4 1 99 0 0 8320 0 97 96 0 0 4
518 470
535 470
535 544
543 544
1 0 80 0 0 4096 0 102 0 0 222 2
399 402
202 402
2 0 94 0 0 4096 0 102 0 0 219 2
399 420
290 420
1 0 79 0 0 4096 0 101 0 0 227 2
482 376
174 376
3 2 100 0 0 4224 0 102 101 0 0 4
445 411
474 411
474 394
482 394
2 0 94 0 0 0 0 103 0 0 219 2
353 361
290 361
1 0 77 0 0 0 0 103 0 0 223 2
353 343
226 343
1 0 78 0 0 4096 0 104 0 0 226 2
478 294
146 294
3 2 101 0 0 8320 0 103 104 0 0 3
408 352
408 312
478 312
2 0 94 0 0 0 0 107 0 0 219 2
374 273
290 273
1 0 82 0 0 0 0 105 0 0 230 2
375 179
116 179
3 2 102 0 0 4224 0 107 106 0 0 4
429 264
464 264
464 230
472 230
0 1 79 0 0 0 0 0 107 227 0 4
174 220
367 220
367 255
374 255
0 2 77 0 0 0 0 0 105 223 0 4
226 260
349 260
349 197
375 197
3 1 103 0 0 4224 0 105 106 0 0 4
421 188
452 188
452 212
472 212
0 1 94 0 0 0 0 0 108 219 0 3
290 109
263 109
263 118
1 0 94 0 0 4224 0 9 0 0 0 2
290 97
290 1209
2 0 81 0 0 4224 0 108 0 0 0 2
263 154
263 1212
1 0 77 0 0 0 0 109 0 0 223 2
202 116
226 116
2 0 80 0 0 4224 0 109 0 0 0 2
202 152
202 1215
1 0 77 0 0 4224 0 10 0 0 0 2
226 95
226 1212
1 0 79 0 0 0 0 110 0 0 227 2
146 113
174 113
1 0 82 0 0 0 0 111 0 0 230 2
85 114
116 114
2 0 78 0 0 4224 0 110 0 0 0 2
146 149
146 1215
1 0 79 0 0 4224 0 11 0 0 0 2
174 94
174 1214
1 0 79 0 0 0 0 11 0 0 0 2
174 94
174 656
2 0 104 0 0 4224 0 111 0 0 0 2
85 150
85 1217
1 0 82 0 0 4224 0 12 0 0 0 2
116 94
116 1216
17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
525 2986 550 3010
533 2994 541 3010
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
568 2727 593 2751
576 2735 584 2751
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
564 2560 589 2584
572 2568 580 2584
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 499 610 523
593 507 601 523
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
518 350 547 374
528 358 536 374
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
529 269 554 293
537 277 545 293
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
527 187 556 211
537 195 545 211
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
576 691 605 715
586 699 594 715
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
581 844 610 868
591 852 599 868
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 1006 614 1030
595 1014 603 1030
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
654 1669 683 1693
664 1677 672 1693
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
591 1995 620 2019
601 2003 609 2019
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
514 2193 539 2217
522 2201 530 2217
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 5 55 29
28 13 44 29
2 a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
239 11 492 35
249 19 481 35
29 Decodificador BCD 7 segmentos
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 37
245 1377 562 1401
255 1385 551 1401
37 Decodificador hexadecimal 7 segmentos
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
614 2375 639 2399
622 2383 630 2399
1 d
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
