CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 489
9437202 0
0
6 Title:
5 Name:
0
0
0
21
9 3-In AND~
219 399 636 0 1 22
0 0
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 6 0
1 U
7762 0 0
2
43728.1 0
0
8 3-In OR~
219 556 553 0 4 22
0 6 5 4 3
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
6723 0 0
2
43728.1 5
0
8 3-In OR~
219 485 470 0 4 22
0 9 8 7 6
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
6871 0 0
2
43728.1 4
0
9 2-In AND~
219 403 481 0 3 22
0 10 11 8
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4198 0 0
2
43728.1 2
0
9 2-In AND~
219 402 530 0 3 22
0 11 12 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
970 0 0
2
43728.1 1
0
9 2-In AND~
219 397 588 0 3 22
0 10 12 5
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
319 0 0
2
43728.1 0
0
13 Logic Switch~
5 290 85 0 1 11
0 25
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3663 0 0
2
43728 0
0
13 Logic Switch~
5 226 83 0 1 11
0 28
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 W
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3512 0 0
2
43728 0
0
13 Logic Switch~
5 174 82 0 1 11
0 26
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7555 0 0
2
43728 0
0
13 Logic Switch~
5 116 82 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-7 -21 7 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9776 0 0
2
43728 0
0
8 2-In OR~
219 495 385 0 3 22
0 26 27 48
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 7 0
1 U
6596 0 0
2
43728.1 1
0
8 2-In OR~
219 412 411 0 3 22
0 24 25 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
6750 0 0
2
43728.1 0
0
6 74266~
219 369 352 0 3 22
0 28 25 30
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9636 0 0
2
43728.1 1
0
8 2-In OR~
219 491 303 0 3 22
0 29 30 49
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 3 0
1 U
5369 0 0
2
43728.1 0
0
8 2-In OR~
219 388 188 0 3 22
0 31 28 33
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8555 0 0
2
43728 6
0
8 2-In OR~
219 485 221 0 3 22
0 33 32 50
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 3 0
1 U
4690 0 0
2
43728 5
0
6 74266~
219 390 264 0 3 22
0 26 25 32
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9145 0 0
2
43728 4
0
9 Inverter~
13 260 136 0 2 22
0 25 34
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
5246 0 0
2
43728 0
0
9 Inverter~
13 199 134 0 2 22
0 28 24
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
9111 0 0
2
43728 0
0
9 Inverter~
13 143 131 0 2 22
0 26 29
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
6717 0 0
2
43728 0
0
9 Inverter~
13 82 132 0 2 22
0 31 35
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3487 0 0
2
43728 0
0
42
3 0 0 0 0 0 0 1 0 0 39 2
375 645
174 645
2 0 0 0 0 0 0 1 0 0 31 2
375 636
290 636
1 0 0 0 0 0 0 1 0 0 34 2
375 627
202 627
2 0 0 0 0 0 0 6 0 0 35 2
373 597
226 597
1 0 0 0 0 0 0 6 0 0 38 2
373 579
146 579
2 0 0 0 0 0 0 5 0 0 32 2
378 539
263 539
1 0 0 0 0 0 0 4 0 0 32 2
379 472
263 472
1 0 0 0 0 0 0 5 0 0 38 2
378 521
146 521
2 0 0 0 0 0 0 4 0 0 35 2
379 490
226 490
3 3 0 0 0 0 0 5 3 0 0 4
423 530
452 530
452 479
472 479
3 2 0 0 0 0 0 4 3 0 0 4
424 481
440 481
440 470
473 470
1 0 0 0 0 0 0 3 0 0 42 2
472 461
116 461
4 3 4 0 0 16 0 1 2 0 0 4
420 636
520 636
520 562
543 562
3 2 5 0 0 0 0 6 2 0 0 4
418 588
495 588
495 553
544 553
4 1 6 0 0 0 0 3 2 0 0 4
518 470
535 470
535 544
543 544
1 0 24 0 0 4096 0 12 0 0 34 2
399 402
202 402
2 0 25 0 0 4096 0 12 0 0 31 2
399 420
290 420
1 0 26 0 0 4096 0 11 0 0 39 2
482 376
174 376
3 2 27 0 0 4224 0 12 11 0 0 4
445 411
474 411
474 394
482 394
2 0 25 0 0 0 0 13 0 0 31 2
353 361
290 361
1 0 28 0 0 4096 0 13 0 0 35 2
353 343
226 343
1 0 29 0 0 4096 0 14 0 0 38 2
478 294
146 294
3 2 30 0 0 8320 0 13 14 0 0 3
408 352
408 312
478 312
2 0 25 0 0 0 0 17 0 0 31 2
374 273
290 273
1 0 31 0 0 4096 0 15 0 0 42 2
375 179
116 179
3 2 32 0 0 4224 0 17 16 0 0 4
429 264
464 264
464 230
472 230
0 1 26 0 0 0 0 0 17 39 0 4
174 220
367 220
367 255
374 255
0 2 28 0 0 0 0 0 15 35 0 4
226 260
349 260
349 197
375 197
3 1 33 0 0 4224 0 15 16 0 0 4
421 188
452 188
452 212
472 212
0 1 25 0 0 0 0 0 18 31 0 3
290 109
263 109
263 118
1 0 25 0 0 4224 0 7 0 0 0 2
290 97
290 670
2 0 34 0 0 4224 0 18 0 0 0 2
263 154
263 675
1 0 28 0 0 0 0 19 0 0 35 2
202 116
226 116
2 0 24 0 0 4224 0 19 0 0 0 2
202 152
202 673
1 0 28 0 0 4224 0 8 0 0 0 2
226 95
226 668
1 0 26 0 0 0 0 20 0 0 39 2
146 113
174 113
1 0 31 0 0 0 0 21 0 0 42 2
85 114
116 114
2 0 29 0 0 4224 0 20 0 0 0 2
146 149
146 670
1 0 26 0 0 4224 0 9 0 0 0 2
174 94
174 670
1 0 26 0 0 0 0 9 0 0 0 2
174 94
174 656
2 0 35 0 0 4224 0 21 0 0 0 2
85 150
85 671
1 0 31 0 0 4224 0 10 0 0 0 2
116 94
116 672
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 499 610 523
593 507 601 523
1 d
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
518 350 547 374
528 358 536 374
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
529 269 554 293
537 277 545 293
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
527 187 556 211
537 195 545 211
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1204 1079 1233 1103
1214 1087 1222 1103
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1299 676 1376 700
1309 684 1365 700
7 SAIDA D
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
