CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
37
13 Logic Switch~
5 290 85 0 1 11
0 27
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Z
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7548 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 226 83 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 W
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8973 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 174 82 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9712 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 116 82 0 1 11
0 15
0
0 0 21360 270
2 0V
-7 -21 7 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4518 0 0
2
5.89908e-315 0
0
7 Ground~
168 813 417 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5596 0 0
2
43728.3 0
0
9 CC 7-Seg~
183 727 380 0 17 19
10 9 8 7 6 5 4 3 38 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
692 0 0
2
43728.3 0
0
8 2-In OR~
219 515 1013 0 3 22
0 15 17 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
6258 0 0
2
43728.3 8
0
8 2-In OR~
219 508 1124 0 3 22
0 19 18 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
5578 0 0
2
43728.3 7
0
8 2-In OR~
219 579 1073 0 3 22
0 20 16 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
8709 0 0
2
43728.3 6
0
9 2-In AND~
219 416 1034 0 3 22
0 10 11 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
9131 0 0
2
43728.3 2
0
9 2-In AND~
219 416 1092 0 3 22
0 12 13 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
3645 0 0
2
43728.3 1
0
9 2-In AND~
219 415 1151 0 3 22
0 10 14 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
7613 0 0
2
43728.3 0
0
8 2-In OR~
219 557 892 0 3 22
0 22 21 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
9467 0 0
2
43728.3 7
0
8 2-In OR~
219 482 930 0 3 22
0 24 23 21
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
3932 0 0
2
43728.3 6
0
8 2-In OR~
219 485 855 0 3 22
0 25 15 22
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
5288 0 0
2
43728.3 5
0
9 2-In AND~
219 409 832 0 3 22
0 12 14 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
4934 0 0
2
43728.3 4
0
9 2-In AND~
219 408 899 0 3 22
0 12 13 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
5987 0 0
2
43728.3 3
0
9 2-In AND~
219 405 958 0 3 22
0 13 14 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
7737 0 0
2
43728.3 2
0
9 2-In AND~
219 553 746 0 3 22
0 26 14 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
4200 0 0
2
43728.3 1
0
8 2-In OR~
219 446 717 0 3 22
0 11 10 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
5780 0 0
2
43728.3 0
0
9 3-In AND~
219 399 636 0 4 22
0 13 27 12 30
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 6 0
1 U
6490 0 0
2
5.89909e-315 0
0
8 3-In OR~
219 556 553 0 4 22
0 32 31 30 6
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
8663 0 0
2
5.89909e-315 5.3568e-315
0
8 3-In OR~
219 485 470 0 4 22
0 15 29 28 32
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
318 0 0
2
5.89909e-315 5.34643e-315
0
9 2-In AND~
219 403 481 0 3 22
0 14 10 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
348 0 0
2
5.89909e-315 5.30499e-315
0
9 2-In AND~
219 402 530 0 3 22
0 11 14 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
8551 0 0
2
5.89909e-315 5.26354e-315
0
9 2-In AND~
219 397 588 0 3 22
0 11 10 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
7295 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 495 385 0 3 22
0 12 33 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
9900 0 0
2
5.89909e-315 5.26354e-315
0
8 2-In OR~
219 412 411 0 3 22
0 13 27 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
8725 0 0
2
5.89909e-315 0
0
6 74266~
219 369 352 0 3 22
0 10 27 34
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
366 0 0
2
5.89909e-315 5.26354e-315
0
8 2-In OR~
219 491 303 0 3 22
0 11 34 8
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
5762 0 0
2
5.89909e-315 0
0
8 2-In OR~
219 388 188 0 3 22
0 15 10 36
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4943 0 0
2
5.89908e-315 5.36716e-315
0
8 2-In OR~
219 485 221 0 3 22
0 36 35 9
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3435 0 0
2
5.89908e-315 5.3568e-315
0
6 74266~
219 390 264 0 3 22
0 12 27 35
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
8705 0 0
2
5.89908e-315 5.34643e-315
0
9 Inverter~
13 260 136 0 2 22
0 27 14
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
4331 0 0
2
5.89908e-315 0
0
9 Inverter~
13 199 134 0 2 22
0 10 13
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U10A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
787 0 0
2
5.89908e-315 0
0
9 Inverter~
13 143 131 0 2 22
0 12 11
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3655 0 0
2
5.89908e-315 0
0
9 Inverter~
13 82 132 0 2 22
0 15 37
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
6682 0 0
2
5.89908e-315 0
0
78
7 3 3 0 0 4224 0 6 9 0 0 3
742 416
742 1073
612 1073
6 3 4 0 0 4224 0 6 13 0 0 3
736 416
736 892
590 892
5 3 5 0 0 4224 0 6 19 0 0 3
730 416
730 746
574 746
4 4 6 0 0 4224 0 6 22 0 0 3
724 416
724 553
589 553
3 3 7 0 0 8320 0 6 27 0 0 5
718 416
718 430
541 430
541 385
528 385
2 3 8 0 0 8320 0 6 30 0 0 5
712 416
712 425
537 425
537 303
524 303
1 3 9 0 0 12416 0 6 32 0 0 5
706 416
706 420
533 420
533 221
518 221
1 9 2 0 0 8320 0 5 6 0 0 4
813 411
813 330
727 330
727 338
1 0 10 0 0 4096 0 10 0 0 71 2
392 1025
226 1025
2 0 11 0 0 4096 0 10 0 0 74 2
392 1043
146 1043
1 0 12 0 0 4096 0 11 0 0 75 2
392 1083
174 1083
2 0 13 0 0 4096 0 11 0 0 70 2
392 1101
202 1101
2 0 14 0 0 4096 0 12 0 0 68 2
391 1160
263 1160
1 0 10 0 0 0 0 12 0 0 71 2
391 1142
226 1142
1 0 15 0 0 4096 0 7 0 0 78 2
502 1004
116 1004
3 2 16 0 0 8320 0 8 9 0 0 4
541 1124
558 1124
558 1082
566 1082
3 2 17 0 0 4224 0 10 7 0 0 4
437 1034
471 1034
471 1022
502 1022
3 2 18 0 0 4224 0 12 8 0 0 4
436 1151
476 1151
476 1133
495 1133
3 1 19 0 0 4224 0 11 8 0 0 4
437 1092
476 1092
476 1115
495 1115
3 1 20 0 0 4224 0 7 9 0 0 3
548 1013
548 1064
566 1064
2 0 14 0 0 0 0 18 0 0 68 2
381 967
263 967
2 0 13 0 0 0 0 17 0 0 70 2
384 908
202 908
1 0 13 0 0 0 0 18 0 0 70 2
381 949
202 949
2 0 14 0 0 0 0 16 0 0 68 2
385 841
263 841
1 0 12 0 0 0 0 16 0 0 75 2
385 823
174 823
2 0 15 0 0 0 0 15 0 0 78 2
472 864
116 864
3 2 21 0 0 8320 0 14 13 0 0 4
515 930
536 930
536 901
544 901
3 1 22 0 0 8320 0 15 13 0 0 4
518 855
536 855
536 883
544 883
3 2 23 0 0 4224 0 18 14 0 0 4
426 958
461 958
461 939
469 939
3 1 24 0 0 4224 0 17 14 0 0 4
429 899
461 899
461 921
469 921
3 1 25 0 0 8320 0 16 15 0 0 3
430 832
430 846
472 846
0 1 12 0 0 0 0 0 17 75 0 2
174 890
384 890
0 2 14 0 0 4096 0 0 19 68 0 4
263 781
513 781
513 755
529 755
3 1 26 0 0 4224 0 20 19 0 0 4
479 717
512 717
512 737
529 737
0 2 10 0 0 4096 0 0 20 71 0 4
226 741
396 741
396 726
433 726
0 1 11 0 0 4096 0 0 20 74 0 4
146 693
396 693
396 708
433 708
3 0 12 0 0 0 0 21 0 0 75 2
375 645
174 645
2 0 27 0 0 4096 0 21 0 0 67 2
375 636
290 636
1 0 13 0 0 0 0 21 0 0 70 2
375 627
202 627
2 0 10 0 0 0 0 26 0 0 71 2
373 597
226 597
1 0 11 0 0 0 0 26 0 0 74 2
373 579
146 579
2 0 14 0 0 0 0 25 0 0 68 2
378 539
263 539
1 0 14 0 0 0 0 24 0 0 68 2
379 472
263 472
1 0 11 0 0 0 0 25 0 0 74 2
378 521
146 521
2 0 10 0 0 0 0 24 0 0 71 2
379 490
226 490
3 3 28 0 0 8320 0 25 23 0 0 4
423 530
452 530
452 479
472 479
3 2 29 0 0 12416 0 24 23 0 0 4
424 481
440 481
440 470
473 470
1 0 15 0 0 0 0 23 0 0 78 2
472 461
116 461
4 3 30 0 0 4224 0 21 22 0 0 4
420 636
520 636
520 562
543 562
3 2 31 0 0 4224 0 26 22 0 0 4
418 588
495 588
495 553
544 553
4 1 32 0 0 8320 0 23 22 0 0 4
518 470
535 470
535 544
543 544
1 0 13 0 0 4096 0 28 0 0 70 2
399 402
202 402
2 0 27 0 0 4096 0 28 0 0 67 2
399 420
290 420
1 0 12 0 0 4096 0 27 0 0 75 2
482 376
174 376
3 2 33 0 0 4224 0 28 27 0 0 4
445 411
474 411
474 394
482 394
2 0 27 0 0 0 0 29 0 0 67 2
353 361
290 361
1 0 10 0 0 0 0 29 0 0 71 2
353 343
226 343
1 0 11 0 0 4096 0 30 0 0 74 2
478 294
146 294
3 2 34 0 0 8320 0 29 30 0 0 3
408 352
408 312
478 312
2 0 27 0 0 0 0 33 0 0 67 2
374 273
290 273
1 0 15 0 0 0 0 31 0 0 78 2
375 179
116 179
3 2 35 0 0 4224 0 33 32 0 0 4
429 264
464 264
464 230
472 230
0 1 12 0 0 0 0 0 33 75 0 4
174 220
367 220
367 255
374 255
0 2 10 0 0 0 0 0 31 71 0 4
226 260
349 260
349 197
375 197
3 1 36 0 0 4224 0 31 32 0 0 4
421 188
452 188
452 212
472 212
0 1 27 0 0 0 0 0 34 67 0 3
290 109
263 109
263 118
1 0 27 0 0 4224 0 1 0 0 0 2
290 97
290 1209
2 0 14 0 0 4224 0 34 0 0 0 2
263 154
263 1212
1 0 10 0 0 0 0 35 0 0 71 2
202 116
226 116
2 0 13 0 0 4224 0 35 0 0 0 2
202 152
202 1215
1 0 10 0 0 4224 0 2 0 0 0 2
226 95
226 1212
1 0 12 0 0 0 0 36 0 0 75 2
146 113
174 113
1 0 15 0 0 0 0 37 0 0 78 2
85 114
116 114
2 0 11 0 0 4224 0 36 0 0 0 2
146 149
146 1215
1 0 12 0 0 4224 0 3 0 0 0 2
174 94
174 1214
1 0 12 0 0 0 0 3 0 0 0 2
174 94
174 656
2 0 37 0 0 4224 0 37 0 0 0 2
85 150
85 1217
1 0 15 0 0 4224 0 4 0 0 0 2
116 94
116 1216
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 1006 614 1030
595 1014 603 1030
1 g
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
581 844 610 868
591 852 599 868
1 f
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
576 691 605 715
586 699 594 715
1 e
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1299 676 1376 700
1309 684 1365 700
7 SAIDA D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1204 1079 1233 1103
1214 1087 1222 1103
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
527 187 556 211
537 195 545 211
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
529 269 554 293
537 277 545 293
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
518 350 547 374
528 358 536 374
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
585 499 610 523
593 507 601 523
1 d
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
