CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 949 95 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-7 -23 7 -15
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43787.9 0
0
6 74LS48
188 311 678 0 14 29
0 2 5 4 3 32 33 12 11 10
9 8 7 6 34
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
3 U13
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
391 0 0
2
5.89916e-315 5.32571e-315
0
7 Ground~
168 243 600 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.89916e-315 5.30499e-315
0
9 CC 7-Seg~
183 434 585 0 17 19
10 6 7 8 9 10 11 12 35 2
1 1 1 1 0 0 1 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3421 0 0
2
5.89916e-315 5.26354e-315
0
7 Ground~
168 434 528 0 1 3
0 2
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8157 0 0
2
5.89916e-315 0
0
5 4082~
219 750 620 0 5 22
0 14 15 16 17 18
0
0 0 624 180
4 4082
-7 -24 21 -16
3 U5A
-13 -28 8 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
5572 0 0
2
5.89916e-315 0
0
5 4071~
219 681 720 0 3 22
0 21 22 3
0
0 0 624 180
4 4071
-7 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
8901 0 0
2
5.89916e-315 0
0
5 4082~
219 746 747 0 5 22
0 14 15 19 17 21
0
0 0 624 180
4 4082
-7 -24 21 -16
3 U4B
-13 -28 8 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
7361 0 0
2
5.89916e-315 0
0
5 4082~
219 745 700 0 5 22
0 14 15 20 17 22
0
0 0 624 180
4 4082
-7 -24 21 -16
3 U4A
-13 -28 8 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
4747 0 0
2
5.89916e-315 0
0
5 4081~
219 751 575 0 3 22
0 20 14 23
0
0 0 624 180
4 4081
-7 -24 21 -16
3 U1B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
972 0 0
2
5.89916e-315 0
0
5 4071~
219 686 597 0 3 22
0 18 23 4
0
0 0 624 180
4 4071
-7 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3472 0 0
2
5.89916e-315 0
0
5 4081~
219 747 496 0 3 22
0 19 14 5
0
0 0 624 180
4 4081
-7 -24 21 -16
3 U1A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9998 0 0
2
5.89916e-315 0
0
2 +V
167 1014 455 0 1 3
0 17
0
0 0 53744 0
2 5V
-8 -22 6 -14
2 V1
-8 -32 6 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
5.89916e-315 0
0
14 Logic Display~
6 669 326 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
43787.9 5
0
14 Logic Display~
6 543 328 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
43787.9 6
0
14 Logic Display~
6 403 331 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
43787.9 7
0
5 4027~
219 613 431 0 7 32
0 36 29 16 29 37 14 26
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U7A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
5616 0 0
2
43787.9 8
0
9 Inverter~
13 981 138 0 2 22
0 15 27
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U8A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
9323 0 0
2
43787.9 9
0
14 Logic Display~
6 193 311 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
43787.9 10
0
7 Pulser~
4 153 395 0 10 12
0 38 39 40 30 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3108 0 0
2
43787.9 11
0
5 4027~
219 344 436 0 7 32
0 41 31 30 31 42 24 20
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
4299 0 0
2
43787.9 12
0
5 4027~
219 488 432 0 7 32
0 43 28 24 28 44 16 19
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
9672 0 0
2
43787.9 13
0
56
3 4 3 0 0 8320 0 7 2 0 0 5
654 720
654 930
275 930
275 669
279 669
3 3 4 0 0 12416 0 11 2 0 0 6
659 597
581 597
581 900
260 900
260 660
279 660
3 2 5 0 0 8320 0 12 2 0 0 6
720 496
547 496
547 860
247 860
247 651
279 651
13 1 6 0 0 8320 0 2 4 0 0 3
343 696
413 696
413 621
12 2 7 0 0 4224 0 2 4 0 0 3
343 687
419 687
419 621
11 3 8 0 0 4224 0 2 4 0 0 3
343 678
425 678
425 621
10 4 9 0 0 4224 0 2 4 0 0 3
343 669
431 669
431 621
9 5 10 0 0 4224 0 2 4 0 0 3
343 660
437 660
437 621
8 6 11 0 0 4224 0 2 4 0 0 3
343 651
443 651
443 621
7 7 12 0 0 4224 0 2 4 0 0 3
343 642
449 642
449 621
1 9 2 0 0 4096 0 5 4 0 0 4
434 536
434 551
434 551
434 543
1 1 2 0 0 4224 0 2 3 0 0 3
279 642
243 642
243 608
0 0 13 0 0 8320 0 0 0 0 0 3
725 499
725 500
719 500
1 0 14 0 0 4096 0 6 0 0 40 2
768 633
902 633
2 0 15 0 0 4096 0 6 0 0 51 2
768 624
949 624
3 0 16 0 0 4096 0 6 0 0 42 2
768 615
852 615
4 0 17 0 0 4096 0 6 0 0 38 2
768 606
1014 606
5 0 18 0 0 4096 0 6 0 0 32 2
723 620
721 620
1 0 14 0 0 4096 0 8 0 0 40 2
764 760
902 760
2 0 15 0 0 4096 0 8 0 0 51 2
764 751
949 751
3 0 19 0 0 4096 0 8 0 0 43 2
764 742
831 742
1 0 14 0 0 4096 0 9 0 0 40 2
763 713
902 713
2 0 15 0 0 4096 0 9 0 0 51 2
763 704
949 704
3 0 20 0 0 4096 0 9 0 0 45 2
763 695
781 695
0 2 15 0 0 0 0 0 8 0 0 3
757 752
757 751
764 751
4 0 17 0 0 4096 0 8 0 0 38 2
764 733
1014 733
4 0 17 0 0 4096 0 9 0 0 38 2
763 686
1014 686
1 5 21 0 0 8320 0 7 8 0 0 3
700 729
700 747
719 747
2 5 22 0 0 8320 0 7 9 0 0 3
700 711
700 700
718 700
1 0 20 0 0 0 0 10 0 0 45 2
769 584
781 584
2 0 14 0 0 0 0 10 0 0 40 2
769 566
902 566
1 0 18 0 0 4224 0 11 0 0 0 4
705 606
721 606
721 620
725 620
2 3 23 0 0 8320 0 11 10 0 0 3
705 588
705 575
724 575
1 0 19 0 0 0 0 12 0 0 43 2
765 505
831 505
2 0 14 0 0 0 0 12 0 0 40 2
765 487
902 487
0 3 16 0 0 0 0 0 17 42 0 2
564 404
589 404
0 3 24 0 0 8192 0 0 22 44 0 3
439 406
439 405
464 405
1 0 17 0 0 4224 0 13 0 0 0 2
1014 464
1014 971
0 0 25 0 0 0 0 0 0 0 0 2
855 962
855 962
6 0 14 0 0 16512 0 17 0 0 0 5
643 413
766 413
766 196
902 196
902 976
0 0 26 0 0 16512 0 0 0 46 0 5
669 386
752 386
752 172
882 172
882 977
6 0 16 0 0 16512 0 22 0 0 0 5
518 414
564 414
564 156
852 156
852 976
1 0 19 0 0 16512 0 15 0 0 0 5
543 346
575 346
575 134
831 134
831 976
6 0 24 0 0 16512 0 21 0 0 0 5
374 418
439 418
439 121
804 121
804 972
0 0 20 0 0 16512 0 0 0 48 0 5
403 361
427 361
427 114
781 114
781 974
7 1 26 0 0 0 0 17 14 0 0 3
637 395
669 395
669 344
7 1 19 0 0 0 0 22 15 0 0 3
512 396
543 396
543 346
7 1 20 0 0 0 0 21 16 0 0 3
368 400
403 400
403 349
1 0 15 0 0 0 0 18 0 0 51 2
984 120
949 120
2 0 27 0 0 12416 0 18 0 0 0 4
984 156
984 495
985 495
985 976
1 0 15 0 0 4224 0 1 0 0 0 2
949 107
949 972
2 4 28 0 0 8320 0 22 22 0 0 4
464 396
454 396
454 414
464 414
2 4 29 0 0 12416 0 17 17 0 0 6
589 395
589 394
578 394
578 412
589 412
589 413
1 0 30 0 0 4096 0 19 0 0 55 2
193 329
193 407
3 4 30 0 0 4224 0 21 20 0 0 5
320 409
193 409
193 407
183 407
183 395
2 4 31 0 0 8320 0 21 21 0 0 4
320 400
313 400
313 418
320 418
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
363 347 392 371
373 355 381 371
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
880 166 917 190
890 174 906 190
2 C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
855 148 884 172
865 156 873 172
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
828 127 865 151
838 135 854 151
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
811 106 840 130
821 114 829 130
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
779 95 816 119
789 103 805 119
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
759 87 788 111
769 95 777 111
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
505 344 534 368
515 352 523 368
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
625 342 654 366
635 350 643 366
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
695 469 734 492
707 479 721 494
2 C+
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
635 569 674 592
647 579 661 594
2 B+
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
628 692 667 715
640 702 654 717
2 A+
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
