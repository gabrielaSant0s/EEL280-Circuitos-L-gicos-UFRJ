CircuitMaker Text
5.6
Probes: 1
U3C_8
Operating Point
0 230 874 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1010 30 100 10
122 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
290 176 1532 489
1083179026 0
0
6 Title:
5 Name:
0
0
0
104
13 Logic Switch~
5 625 1318 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 B8
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7643 0 0
2
43723.9 1
0
13 Logic Switch~
5 625 1256 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 A8
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3236 0 0
2
43723.9 0
0
13 Logic Switch~
5 86 1268 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 A1
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3903 0 0
2
43723.9 1
0
13 Logic Switch~
5 86 1330 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 B1
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3968 0 0
2
43723.9 0
0
13 Logic Switch~
5 688 1088 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
3 E12
-33 -15 -12 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3106 0 0
2
43723.9 0
0
13 Logic Switch~
5 692 1040 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 D8
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3223 0 0
2
43723.9 0
0
13 Logic Switch~
5 691 890 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-33 -3 -19 5
2 A7
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6341 0 0
2
43723.9 2
0
13 Logic Switch~
5 691 949 0 1 11
0 25
0
0 0 21344 0
2 0V
-28 0 -14 8
2 B7
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4627 0 0
2
43723.9 1
0
13 Logic Switch~
5 693 995 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 C7
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6952 0 0
2
43723.9 0
0
13 Logic Switch~
5 687 732 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 C6
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3974 0 0
2
43723.8 2
0
13 Logic Switch~
5 685 686 0 1 11
0 33
0
0 0 21344 0
2 0V
-28 0 -14 8
2 B6
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4630 0 0
2
43723.8 1
0
13 Logic Switch~
5 686 653 0 1 11
0 34
0
0 0 21344 0
2 0V
-33 -3 -19 5
2 A6
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5705 0 0
2
43723.8 0
0
13 Logic Switch~
5 686 496 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 D5
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8423 0 0
2
43723.8 0
0
13 Logic Switch~
5 686 449 0 1 11
0 45
0
0 0 21344 0
2 0V
-29 -1 -15 7
2 C5
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6486 0 0
2
43723.7 2
0
13 Logic Switch~
5 690 387 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-28 0 -14 8
2 B5
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3367 0 0
2
43723.7 1
0
13 Logic Switch~
5 686 329 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-33 -3 -19 5
2 A5
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7389 0 0
2
43723.7 0
0
13 Logic Switch~
5 706 131 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-33 -3 -19 5
2 A4
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6782 0 0
2
43723.7 2
0
13 Logic Switch~
5 705 164 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-28 0 -14 8
2 B4
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5728 0 0
2
43723.7 1
0
13 Logic Switch~
5 707 210 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-29 -1 -15 7
2 C4
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6119 0 0
2
43723.7 0
0
13 Logic Switch~
5 65 1046 0 1 11
0 57
0
0 0 21360 0
2 0V
-29 -1 -15 7
2 E5
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3241 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 65 1003 0 1 11
0 56
0
0 0 21360 0
2 0V
-29 -1 -15 7
2 D4
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3835 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 63 949 0 1 11
0 60
0
0 0 21360 0
2 0V
-29 -1 -15 7
2 C3
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7478 0 0
2
5.89908e-315 5.30499e-315
0
13 Logic Switch~
5 61 898 0 1 11
0 61
0
0 0 21360 0
2 0V
-28 0 -14 8
2 B3
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3979 0 0
2
5.89908e-315 5.26354e-315
0
13 Logic Switch~
5 62 865 0 1 11
0 64
0
0 0 21360 0
2 0V
-33 -3 -19 5
2 A3
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6285 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 84 481 0 10 11
0 69 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 -1 -15 7
2 D2
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4935 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 77 273 0 1 11
0 71
0
0 0 21360 0
2 0V
-33 -3 -19 5
2 A2
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7650 0 0
2
5.89908e-315 5.30499e-315
0
13 Logic Switch~
5 76 306 0 1 11
0 74
0
0 0 21360 0
2 0V
-28 0 -14 8
2 B2
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9836 0 0
2
5.89908e-315 5.26354e-315
0
13 Logic Switch~
5 78 352 0 10 11
0 73 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 -1 -15 7
2 C2
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3988 0 0
2
5.89908e-315 0
0
13 Logic Switch~
5 81 186 0 10 11
0 76 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 -1 -15 7
2 C1
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
492 0 0
2
5.89908e-315 5.32571e-315
0
13 Logic Switch~
5 79 140 0 10 11
0 75 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-28 0 -14 8
2 B1
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5338 0 0
2
5.89908e-315 5.30499e-315
0
13 Logic Switch~
5 80 107 0 10 11
0 81 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-33 -3 -19 5
2 A1
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8324 0 0
2
5.89908e-315 5.26354e-315
0
13 Logic Switch~
5 78 639 0 1 11
0 87
0
0 0 21360 0
2 0V
-33 -3 -19 5
2 A3
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9550 0 0
2
5.89908e-315 5.3568e-315
0
13 Logic Switch~
5 77 672 0 1 11
0 85
0
0 0 21360 0
2 0V
-28 0 -14 8
2 B3
-28 -14 -14 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6380 0 0
2
5.89908e-315 5.34643e-315
0
13 Logic Switch~
5 79 718 0 10 11
0 86 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 -1 -15 7
2 C3
-30 -15 -16 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7942 0 0
2
5.89908e-315 5.32571e-315
0
7 Ground~
168 1083 1338 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
789 0 0
2
43723.9 1
0
4 LED~
171 1083 1301 0 2 2
10 3 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
9884 0 0
2
43723.9 0
0
5 4011~
219 1020 1269 0 3 22
0 4 4 3
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U23B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 23 0
1 U
6253 0 0
2
43723.9 0
0
5 4011~
219 822 1306 0 3 22
0 7 8 5
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U23A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 23 0
1 U
7409 0 0
2
43723.9 0
0
5 4011~
219 715 1309 0 3 22
0 8 8 9
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U22D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 22 0
1 U
3540 0 0
2
43723.9 0
0
5 4011~
219 717 1246 0 3 22
0 7 7 10
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U22C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 22 0
1 U
3103 0 0
2
43723.9 0
0
5 4011~
219 926 1278 0 3 22
0 6 5 4
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U22B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 22 0
1 U
3548 0 0
2
43723.9 0
0
5 4011~
219 821 1256 0 3 22
0 10 9 6
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U22A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 22 0
1 U
9961 0 0
2
43723.9 0
0
4 LED~
171 351 1321 0 2 2
10 12 11
0
0 0 880 0
4 LED1
17 1 45 9
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8521 0 0
2
43723.9 6
0
2 +V
167 352 1243 0 1 3
0 13
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5296 0 0
2
43723.9 5
0
5 4001~
219 257 1290 0 3 22
0 15 14 11
0
0 0 608 0
4 4001
-14 -24 14 -16
4 U12C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 12 0
1 U
5398 0 0
2
43723.9 4
0
9 2-In AND~
219 173 1321 0 3 22
0 17 16 14
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U20B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
7935 0 0
2
43723.9 3
0
9 2-In AND~
219 172 1278 0 3 22
0 17 16 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U20A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
356 0 0
2
43723.9 2
0
4 LED~
171 1100 1005 0 2 2
10 18 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D12
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4629 0 0
2
43723.9 1
0
7 Ground~
168 1100 1042 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
538 0 0
2
43723.9 0
0
5 7422~
219 1036 973 0 5 22
0 22 20 21 19 18
0
0 0 608 0
6 74LS22
-21 -28 21 -20
4 U21A
-15 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 20 0
1 U
5713 0 0
2
43723.9 0
0
5 4011~
219 898 967 0 3 22
0 24 23 21
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U19D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 19 0
1 U
6618 0 0
2
43723.9 0
0
5 4011~
219 895 902 0 3 22
0 26 25 22
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U19C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 19 0
1 U
3714 0 0
2
43723.9 0
0
5 4011~
219 785 1097 0 3 22
0 27 27 19
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U19B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 19 0
1 U
9116 0 0
2
43723.9 0
0
5 4011~
219 787 1006 0 3 22
0 28 28 23
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U19A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 19 0
1 U
7960 0 0
2
43723.9 0
0
5 4011~
219 791 958 0 3 22
0 25 25 24
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 18 0
1 U
3886 0 0
2
43723.9 0
0
5 4011~
219 790 879 0 3 22
0 29 29 26
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 18 0
1 U
3299 0 0
2
43723.9 0
0
7 Ground~
168 969 746 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9107 0 0
2
43723.8 1
0
4 LED~
171 969 709 0 2 2
10 30 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D11
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
6556 0 0
2
43723.8 0
0
10 3-In NAND~
219 904 677 0 4 22
0 32 31 35 30
0
0 0 608 0
5 74F10
-18 -28 17 -20
4 U17B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 17 0
1 U
3205 0 0
2
43723.8 0
0
5 4011~
219 794 693 0 3 22
0 33 33 31
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 18 0
1 U
7255 0 0
2
43723.8 0
0
5 4011~
219 792 644 0 3 22
0 34 34 32
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 18 0
1 U
8613 0 0
2
43723.8 0
0
4 LED~
171 1115 395 0 2 2
10 36 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D10
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
7832 0 0
2
43723.8 1
0
7 Ground~
168 1115 432 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8937 0 0
2
43723.8 0
0
10 3-In NAND~
219 908 486 0 4 22
0 39 38 37 42
0
0 0 608 0
5 74F10
-18 -28 17 -20
4 U17A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 17 0
1 U
556 0 0
2
43723.7 0
0
10 3-In NAND~
219 908 420 0 4 22
0 41 38 40 43
0
0 0 608 0
5 74F10
-18 -28 17 -20
4 U15C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 15 0
1 U
6981 0 0
2
43723.7 0
0
10 3-In NAND~
219 1051 363 0 4 22
0 44 43 42 36
0
0 0 608 0
5 74F10
-18 -28 17 -20
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 15 0
1 U
8701 0 0
2
43723.7 0
0
10 3-In NAND~
219 909 344 0 4 22
0 39 38 40 44
0
0 0 608 0
5 74F10
-18 -28 17 -20
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 15 0
1 U
5540 0 0
2
43723.7 0
0
5 4011~
219 762 448 0 3 22
0 45 45 40
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 14 0
1 U
8365 0 0
2
43723.7 0
0
5 4011~
219 762 387 0 3 22
0 46 46 38
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 14 0
1 U
5209 0 0
2
43723.7 0
0
5 4011~
219 764 320 0 3 22
0 41 41 39
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 14 0
1 U
3297 0 0
2
43723.7 0
0
5 4011~
219 955 165 0 3 22
0 48 48 47
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 14 0
1 U
9904 0 0
2
43723.7 0
0
7 Ground~
168 1018 234 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6918 0 0
2
43723.7 1
0
4 LED~
171 1020 174 0 2 2
10 47 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D9
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
7751 0 0
2
43723.7 0
0
5 4023~
219 852 163 0 4 22
0 49 51 50 48
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U16A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 16 0
1 U
9907 0 0
2
43723.7 0
0
4 LED~
171 403 689 0 2 2
10 53 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
6628 0 0
2
43723.6 0
0
4 LED~
171 491 375 0 2 2
10 54 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
4914 0 0
2
43723.6 0
0
4 LED~
171 466 189 0 2 2
10 52 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
635 0 0
2
43723.6 0
0
4 LED~
171 439 926 0 2 2
10 63 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3606 0 0
2
5.89908e-315 0
0
12 4-In AND:DM~
219 317 902 0 5 22
0 59 58 56 55 63
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 10 0
1 U
8769 0 0
2
5.89908e-315 0
0
11 2-In OR:DM~
219 203 936 0 3 22
0 61 60 58
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
3887 0 0
2
5.89908e-315 0
0
9 Inverter~
13 153 1046 0 2 22
0 57 55
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9B
-11 12 10 20
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
4266 0 0
2
5.89908e-315 0
0
9 Inverter~
13 114 866 0 2 22
0 64 62
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
3389 0 0
2
5.89908e-315 0
0
10 2-In NAND~
219 196 875 0 3 22
0 62 61 59
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8108 0 0
2
5.89908e-315 0
0
7 Ground~
168 439 963 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3301 0 0
2
5.89908e-315 0
0
7 Ground~
168 490 409 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3739 0 0
2
5.89908e-315 5.26354e-315
0
8 3-In OR~
219 406 357 0 4 22
0 72 67 66 54
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
4610 0 0
2
5.89908e-315 0
0
9 3-In AND~
219 272 471 0 4 22
0 65 68 69 66
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 7 0
1 U
7104 0 0
2
5.89908e-315 0
0
9 3-In AND~
219 269 384 0 4 22
0 71 68 70 67
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 5 0
1 U
5233 0 0
2
5.89908e-315 0
0
9 3-In AND~
219 269 284 0 4 22
0 65 68 70 72
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 5 0
1 U
345 0 0
2
5.89908e-315 0
0
9 Inverter~
13 150 352 0 2 22
0 73 70
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6D
-9 12 12 20
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
4311 0 0
2
5.89908e-315 0
0
9 Inverter~
13 150 306 0 2 22
0 74 68
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6C
-9 12 12 20
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
3959 0 0
2
5.89908e-315 0
0
9 Inverter~
13 150 274 0 2 22
0 71 65
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6B
-9 12 12 20
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
9550 0 0
2
5.89908e-315 0
0
9 Inverter~
13 141 140 0 2 22
0 75 79
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-9 12 12 20
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
4183 0 0
2
5.89908e-315 0
0
9 3-In AND~
219 379 178 0 4 22
0 77 75 76 52
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
7662 0 0
2
5.89908e-315 0
0
9 Inverter~
13 262 118 0 2 22
0 78 77
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
6373 0 0
2
5.89908e-315 0
0
8 2-In OR~
219 193 117 0 3 22
0 80 79 78
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
76 0 0
2
5.89908e-315 0
0
9 Inverter~
13 123 107 0 2 22
0 81 80
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
4168 0 0
2
5.89908e-315 0
0
7 Ground~
168 466 222 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9490 0 0
2
5.89908e-315 0
0
9 2-In NOR~
219 204 649 0 3 22
0 87 85 88
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 512 4 4 1 0
1 U
3202 0 0
2
5.89908e-315 5.38788e-315
0
9 2-In NOR~
219 205 710 0 3 22
0 85 84 82
0
0 0 624 0
4 7428
-14 -24 14 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5212 0 0
2
5.89908e-315 5.37752e-315
0
9 Inverter~
13 133 719 0 2 22
0 86 84
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-10 15 11 23
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
5341 0 0
2
5.89908e-315 5.36716e-315
0
10 2-In NAND~
219 321 675 0 3 22
0 83 82 53
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3516 0 0
2
5.89908e-315 5.30499e-315
0
7 Ground~
168 404 723 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6823 0 0
2
5.89908e-315 5.26354e-315
0
9 Resistor~
219 351 1279 0 4 5
0 12 13 0 1
0
0 0 864 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3532 0 0
2
43723.9 7
0
126
3 1 3 0 0 4240 0 37 36 0 0 3
1047 1269
1083 1269
1083 1291
2 1 2 0 0 4112 0 36 35 0 0 2
1083 1311
1083 1332
1 0 4 0 0 4096 0 37 0 0 4 3
996 1260
967 1260
967 1278
3 2 4 0 0 4224 0 41 37 0 0 2
953 1278
996 1278
3 2 5 0 0 4224 0 38 41 0 0 4
849 1306
879 1306
879 1287
902 1287
3 1 6 0 0 4224 0 42 41 0 0 4
848 1256
879 1256
879 1269
902 1269
0 1 7 0 0 16512 0 0 38 14 0 7
653 1255
653 1215
573 1215
573 1361
786 1361
786 1297
798 1297
0 2 8 0 0 8320 0 0 38 12 0 5
647 1318
647 1338
774 1338
774 1315
798 1315
3 2 9 0 0 8320 0 39 42 0 0 4
742 1309
757 1309
757 1265
797 1265
3 1 10 0 0 12416 0 40 42 0 0 4
744 1246
759 1246
759 1247
797 1247
1 0 8 0 0 0 0 39 0 0 12 3
691 1300
665 1300
665 1318
1 2 8 0 0 128 0 1 39 0 0 2
637 1318
691 1318
1 0 7 0 0 0 0 40 0 0 14 3
693 1237
665 1237
665 1255
1 2 7 0 0 128 0 2 40 0 0 3
637 1256
637 1255
693 1255
2 3 11 0 0 4224 0 43 45 0 0 3
351 1331
296 1331
296 1290
1 1 12 0 0 4224 0 104 43 0 0 2
351 1297
351 1311
1 2 13 0 0 8320 0 44 104 0 0 3
352 1252
351 1252
351 1261
3 2 14 0 0 4224 0 46 45 0 0 4
194 1321
221 1321
221 1299
244 1299
3 1 15 0 0 8320 0 47 45 0 0 3
193 1278
193 1281
244 1281
2 0 16 0 0 8192 0 47 0 0 22 3
148 1287
129 1287
129 1330
1 0 17 0 0 8192 0 46 0 0 23 3
149 1312
111 1312
111 1269
1 2 16 0 0 4224 0 4 46 0 0 2
98 1330
149 1330
1 1 17 0 0 8320 0 3 47 0 0 3
98 1268
98 1269
148 1269
5 1 18 0 0 4224 0 50 48 0 0 3
1063 973
1100 973
1100 995
2 1 2 0 0 0 0 48 49 0 0 2
1100 1015
1100 1036
3 4 19 0 0 4224 0 53 50 0 0 4
812 1097
984 1097
984 991
1012 991
1 2 20 0 0 4224 0 6 50 0 0 4
704 1040
933 1040
933 979
1012 979
3 3 21 0 0 4224 0 51 50 0 0 2
925 967
1012 967
3 1 22 0 0 4224 0 52 50 0 0 4
922 902
984 902
984 955
1012 955
3 2 23 0 0 4224 0 54 51 0 0 4
814 1006
847 1006
847 976
874 976
3 1 24 0 0 4224 0 55 51 0 0 2
818 958
874 958
0 2 25 0 0 8320 0 0 52 39 0 3
713 949
713 911
871 911
3 1 26 0 0 4224 0 56 52 0 0 4
817 879
847 879
847 893
871 893
2 0 27 0 0 4096 0 53 0 0 35 3
761 1106
739 1106
739 1088
1 1 27 0 0 4224 0 5 53 0 0 2
700 1088
761 1088
2 0 28 0 0 4096 0 54 0 0 37 3
763 1015
740 1015
740 997
1 1 28 0 0 8320 0 9 54 0 0 3
705 995
705 997
763 997
2 0 25 0 0 0 0 55 0 0 39 3
767 967
739 967
739 949
1 1 25 0 0 128 0 8 55 0 0 2
703 949
767 949
1 0 29 0 0 4096 0 56 0 0 41 3
766 870
739 870
739 888
1 2 29 0 0 8320 0 7 56 0 0 3
703 890
703 888
766 888
4 1 30 0 0 4224 0 59 58 0 0 3
931 677
969 677
969 699
2 1 2 0 0 0 0 58 57 0 0 2
969 719
969 740
3 2 31 0 0 12416 0 60 59 0 0 4
821 693
846 693
846 677
880 677
3 1 32 0 0 12416 0 61 59 0 0 4
819 644
846 644
846 668
880 668
2 0 33 0 0 4096 0 60 0 0 47 3
770 702
735 702
735 684
1 1 33 0 0 8320 0 11 60 0 0 3
697 686
697 684
770 684
1 0 34 0 0 4096 0 61 0 0 49 3
768 635
736 635
736 653
1 2 34 0 0 4224 0 12 61 0 0 2
698 653
768 653
1 3 35 0 0 8320 0 10 59 0 0 5
699 732
699 733
861 733
861 686
880 686
4 1 36 0 0 12416 0 66 62 0 0 5
1078 363
1077 363
1077 363
1115 363
1115 385
2 1 2 0 0 0 0 62 63 0 0 2
1115 405
1115 426
3 1 37 0 0 8320 0 64 13 0 0 3
884 495
884 496
698 496
0 2 38 0 0 4096 0 0 64 57 0 3
833 420
833 486
884 486
1 0 39 0 0 4224 0 64 0 0 64 5
884 477
638 477
638 282
811 282
811 320
3 0 40 0 0 4096 0 65 0 0 62 3
884 429
810 429
810 448
0 2 38 0 0 8320 0 0 65 63 0 3
809 387
809 420
884 420
0 1 41 0 0 8320 0 0 65 70 0 3
711 329
711 411
884 411
4 3 42 0 0 8320 0 64 66 0 0 4
935 486
1003 486
1003 372
1027 372
4 2 43 0 0 8320 0 65 66 0 0 4
935 420
986 420
986 363
1027 363
4 1 44 0 0 4224 0 67 66 0 0 4
936 344
987 344
987 354
1027 354
3 3 40 0 0 8320 0 68 67 0 0 4
789 448
868 448
868 353
885 353
3 2 38 0 0 128 0 69 67 0 0 4
789 387
846 387
846 344
885 344
3 1 39 0 0 128 0 70 67 0 0 4
791 320
847 320
847 335
885 335
1 0 45 0 0 8192 0 68 0 0 66 3
738 439
723 439
723 457
2 1 45 0 0 4224 0 68 14 0 0 3
738 457
698 457
698 449
1 0 46 0 0 8192 0 69 0 0 68 3
738 378
723 378
723 396
2 1 46 0 0 4224 0 69 15 0 0 3
738 396
702 396
702 387
1 0 41 0 0 0 0 70 0 0 70 3
740 311
723 311
723 329
1 2 41 0 0 128 0 16 70 0 0 2
698 329
740 329
3 1 47 0 0 8320 0 71 73 0 0 3
982 165
982 164
1020 164
2 0 48 0 0 4224 0 71 0 0 73 3
931 174
888 174
888 163
4 1 48 0 0 128 0 74 71 0 0 4
879 163
902 163
902 156
931 156
2 1 2 0 0 4224 0 73 72 0 0 3
1020 184
1020 228
1018 228
0 1 49 0 0 4224 0 0 74 78 0 4
728 131
785 131
785 154
828 154
1 3 50 0 0 4224 0 19 74 0 0 4
719 210
785 210
785 172
828 172
1 2 51 0 0 4224 0 18 74 0 0 3
717 164
828 164
828 163
1 1 49 0 0 128 0 17 0 0 0 2
718 131
734 131
4 1 52 0 0 8320 0 94 77 0 0 3
400 178
400 179
466 179
2 1 2 0 0 128 0 75 103 0 0 3
403 699
404 699
404 717
3 1 53 0 0 4224 0 102 75 0 0 4
348 675
404 675
404 679
403 679
2 1 2 0 0 128 0 76 85 0 0 3
491 385
491 403
490 403
4 1 54 0 0 4224 0 86 76 0 0 4
439 357
492 357
492 365
491 365
2 1 2 0 0 0 0 77 98 0 0 2
466 199
466 216
2 1 2 0 0 128 0 78 84 0 0 2
439 936
439 957
2 4 55 0 0 8320 0 81 79 0 0 4
174 1046
281 1046
281 916
296 916
1 3 56 0 0 4224 0 21 79 0 0 4
77 1003
264 1003
264 907
299 907
1 1 57 0 0 4224 0 20 81 0 0 2
77 1046
138 1046
2 3 58 0 0 4224 0 79 80 0 0 4
299 898
243 898
243 936
230 936
3 1 59 0 0 12416 0 83 79 0 0 6
223 875
243 875
243 883
282 883
282 889
296 889
1 2 60 0 0 8320 0 22 80 0 0 3
75 949
75 945
173 945
0 1 61 0 0 8320 0 0 80 95 0 3
88 898
88 927
173 927
2 1 62 0 0 4224 0 82 83 0 0 2
135 866
172 866
5 1 63 0 0 4224 0 79 78 0 0 3
356 902
439 902
439 916
2 1 61 0 0 0 0 83 23 0 0 4
172 884
103 884
103 898
73 898
1 1 64 0 0 8320 0 24 82 0 0 3
74 865
74 866
99 866
1 0 65 0 0 8320 0 87 0 0 108 3
248 462
180 462
180 275
4 3 66 0 0 8320 0 87 86 0 0 4
293 471
356 471
356 366
393 366
4 2 67 0 0 12416 0 88 86 0 0 4
290 384
329 384
329 357
394 357
2 0 68 0 0 4096 0 88 0 0 101 2
245 384
193 384
2 0 68 0 0 8320 0 87 0 0 107 3
248 471
193 471
193 306
3 1 69 0 0 8320 0 87 25 0 0 3
248 480
248 481
96 481
3 0 70 0 0 8192 0 88 0 0 106 3
245 393
220 393
220 352
1 0 71 0 0 4224 0 88 0 0 111 3
245 375
112 375
112 274
4 1 72 0 0 4224 0 89 86 0 0 4
290 284
355 284
355 348
393 348
2 3 70 0 0 4224 0 90 89 0 0 4
171 352
232 352
232 293
245 293
2 2 68 0 0 0 0 91 89 0 0 4
171 306
212 306
212 284
245 284
2 1 65 0 0 0 0 92 89 0 0 3
171 274
171 275
245 275
1 1 73 0 0 4224 0 28 90 0 0 2
90 352
135 352
1 1 74 0 0 4224 0 27 91 0 0 2
88 306
135 306
1 1 71 0 0 0 0 26 92 0 0 3
89 273
89 274
135 274
2 0 75 0 0 4224 0 94 0 0 117 3
355 178
100 178
100 140
3 1 76 0 0 4224 0 94 29 0 0 3
355 187
93 187
93 186
2 1 77 0 0 12416 0 95 94 0 0 4
283 118
296 118
296 169
355 169
3 1 78 0 0 8320 0 96 95 0 0 3
226 117
226 118
247 118
2 2 79 0 0 8320 0 93 96 0 0 3
162 140
162 126
180 126
1 1 75 0 0 0 0 30 93 0 0 2
91 140
126 140
2 1 80 0 0 8320 0 97 96 0 0 3
144 107
144 108
180 108
1 1 81 0 0 4224 0 31 97 0 0 2
92 107
108 107
3 2 82 0 0 4224 0 100 102 0 0 4
244 710
277 710
277 684
297 684
0 1 83 0 0 4224 0 0 102 0 0 4
246 649
278 649
278 666
297 666
2 2 84 0 0 4224 0 101 100 0 0 2
154 719
192 719
1 0 85 0 0 4224 0 100 0 0 125 3
192 701
104 701
104 672
1 1 86 0 0 8320 0 34 101 0 0 3
91 718
91 719
118 719
2 1 85 0 0 0 0 99 33 0 0 4
191 658
119 658
119 672
89 672
1 1 87 0 0 8320 0 32 99 0 0 3
90 639
90 640
191 640
17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 55
648 1159 989 1203
658 1167 978 1199
55 CIRCUITO REDUZIDO APENAS COM PORTAS NAND 
- PAGINA 18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
125 1158 402 1182
135 1166 391 1182
32 FUNCAO COMBINACIONAL - PAGINA 18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 55
698 798 1039 842
708 806 1028 838
55 CIRCUITO REDUZIDO APENAS COM PORTAS NAND 
- PAGINA 17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 55
713 557 1054 601
723 565 1043 597
55 CIRCUITO REDUZIDO APENAS COM PORTAS NAND 
- PAGINA 16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
626 68 663 92
636 76 652 92
2 1)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
580 251 617 275
590 259 606 275
2 2)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 55
728 30 1069 74
738 38 1058 70
55 CIRCUITO REDUZIDO APENAS COM PORTAS NAND 
- PAGINA 15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 142
9 523 1166 547
19 531 1155 547
142 #---------------------------------------------------------------------------------------------------------------------------------------------
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
180 559 457 583
190 567 446 583
32 FUNCAO COMBINACIONAL - PAGINA 16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
359 637 388 661
369 645 377 661
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
192 31 469 55
202 39 458 55
32 FUNCAO COMBINACIONAL - PAGINA 15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
9 58 46 82
19 66 35 82
2 1)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
420 140 449 164
430 148 438 164
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-2 230 35 254
8 238 24 254
2 2)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
445 323 474 347
455 331 463 347
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
178 803 455 827
188 811 444 827
32 FUNCAO COMBINACIONAL - PAGINA 17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
356 869 385 893
366 877 374 893
1 X
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
