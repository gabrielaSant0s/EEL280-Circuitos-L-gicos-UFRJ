CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
43
13 Logic Switch~
5 1052 429 0 1 11
0 28
0
0 0 21360 270
2 0V
-7 -23 7 -15
2 X1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6866 0 0
2
5.89916e-315 0
0
13 Logic Switch~
5 949 95 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-7 -23 7 -15
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7670 0 0
2
5.89916e-315 0
0
6 74LS48
188 1105 503 0 14 29
0 28 17 16 12 47 48 3 4 5
6 7 8 9 49
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
951 0 0
2
43786.7 0
0
14 Logic Display~
6 518 257 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9536 0 0
2
5.89916e-315 0
0
14 Logic Display~
6 258 489 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5495 0 0
2
5.89916e-315 0
0
14 Logic Display~
6 681 1081 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8152 0 0
2
5.89916e-315 5.3568e-315
0
10 2-In NAND~
219 757 1103 0 3 22
0 50 51 20
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U1D
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 1 0
1 U
6223 0 0
2
5.89916e-315 5.34643e-315
0
14 Logic Display~
6 689 1181 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5441 0 0
2
5.89916e-315 5.32571e-315
0
10 2-In NAND~
219 844 1172 0 3 22
0 52 53 23
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U1C
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 1 0
1 U
3189 0 0
2
5.89916e-315 5.30499e-315
0
10 2-In NAND~
219 840 1240 0 3 22
0 54 55 22
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U1B
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 1 0
1 U
8460 0 0
2
5.89916e-315 5.26354e-315
0
10 2-In NAND~
219 766 1203 0 3 22
0 22 23 21
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U1A
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5179 0 0
2
5.89916e-315 0
0
14 Logic Display~
6 420 1072 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3593 0 0
2
5.89916e-315 5.30499e-315
0
10 2-In NAND~
219 570 1061 0 3 22
0 56 57 25
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U6C
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 6 0
1 U
3928 0 0
2
5.89916e-315 5.26354e-315
0
10 2-In NAND~
219 496 1094 0 3 22
0 58 25 24
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U6B
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 6 0
1 U
363 0 0
2
5.89916e-315 0
0
10 2-In NAND~
219 712 270 0 3 22
0 16 26 30
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U6D
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
8132 0 0
2
5.89916e-315 5.32571e-315
0
10 2-In NAND~
219 708 216 0 3 22
0 17 27 31
0
0 0 624 180
6 74LS37
-14 -24 28 -16
4 U10A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
65 0 0
2
5.89916e-315 5.30499e-315
0
10 2-In NAND~
219 713 332 0 3 22
0 12 26 29
0
0 0 624 180
6 74LS37
-14 -24 28 -16
4 U10B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
6609 0 0
2
5.89916e-315 5.26354e-315
0
10 4-In NAND~
219 614 275 0 5 22
0 29 29 30 31 59
0
0 0 624 180
6 74LS20
-21 -28 21 -20
3 U4B
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 512 2 2 4 0
1 U
8995 0 0
2
5.89916e-315 0
0
10 2-In NAND~
219 274 946 0 3 22
0 60 61 37
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U3A
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 3 0
1 U
3918 0 0
2
5.89916e-315 5.38788e-315
0
10 2-In NAND~
219 275 994 0 3 22
0 62 63 36
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U3B
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 3 0
1 U
7519 0 0
2
5.89916e-315 5.37752e-315
0
10 2-In NAND~
219 276 1043 0 3 22
0 64 65 35
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U3C
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 3 0
1 U
377 0 0
2
5.89916e-315 5.36716e-315
0
10 4-In NAND~
219 191 984 0 5 22
0 35 35 36 37 38
0
0 0 624 180
6 74LS20
-21 -28 21 -20
3 U4A
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
8816 0 0
2
5.89916e-315 5.3568e-315
0
14 Logic Display~
6 116 962 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3877 0 0
2
5.89916e-315 5.34643e-315
0
10 2-In NAND~
219 265 1164 0 3 22
0 66 67 33
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U3D
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 3 0
1 U
926 0 0
2
5.89916e-315 5.32571e-315
0
10 2-In XNOR~
219 263 1091 0 3 22
0 68 69 34
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U5A
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 1 5 0
1 U
7262 0 0
2
5.89916e-315 5.30499e-315
0
10 2-In NAND~
219 188 1122 0 3 22
0 33 34 32
0
0 0 624 180
6 74LS37
-14 -24 28 -16
3 U6A
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5267 0 0
2
5.89916e-315 5.26354e-315
0
14 Logic Display~
6 114 1100 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8838 0 0
2
5.89916e-315 0
0
10 2-In NAND~
219 609 774 0 3 22
0 12 17 42
0
0 0 624 180
6 74LS37
-14 -24 28 -16
4 U12A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
7159 0 0
2
5.89916e-315 5.34643e-315
0
10 2-In NAND~
219 612 688 0 3 22
0 17 27 41
0
0 0 624 180
6 74LS37
-14 -24 28 -16
4 U10D
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
5812 0 0
2
5.89916e-315 5.32571e-315
0
10 2-In NAND~
219 610 731 0 3 22
0 12 27 40
0
0 0 624 180
6 74LS37
-14 -24 28 -16
4 U10C
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
331 0 0
2
5.89916e-315 5.30499e-315
0
10 4-In NAND~
219 614 639 0 5 22
0 11 16 26 26 39
0
0 0 624 180
6 74LS20
-21 -28 21 -20
4 U11B
-11 -28 17 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 10 0
1 U
9604 0 0
2
5.89916e-315 5.26354e-315
0
10 4-In NAND~
219 504 714 0 5 22
0 42 40 41 39 13
0
0 0 624 180
6 74LS20
-21 -28 21 -20
4 U11A
-11 -28 17 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 10 0
1 U
7518 0 0
2
5.89916e-315 0
0
9 Inverter~
13 981 138 0 2 22
0 26 27
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U8A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
4832 0 0
2
5.89916e-315 5.26354e-315
0
10 2-In NAND~
219 351 504 0 3 22
0 44 27 70
0
0 0 624 180
6 74LS37
-14 -24 28 -16
4 U12C
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 11 0
1 U
6798 0 0
2
5.89916e-315 5.26354e-315
0
10 2-In NAND~
219 433 536 0 3 22
0 43 27 44
0
0 0 624 180
6 74LS37
-14 -24 28 -16
4 U12B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3336 0 0
2
5.89916e-315 0
0
7 Ground~
168 1232 327 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8370 0 0
2
5.89916e-315 0
0
9 CC 7-Seg~
183 1232 398 0 17 19
10 9 8 7 6 5 4 3 71 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3910 0 0
2
5.89916e-315 5.26354e-315
0
14 Logic Display~
6 91 215 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
316 0 0
2
5.89916e-315 0
0
14 Logic Display~
6 193 311 0 1 2
10 46
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
536 0 0
2
5.89916e-315 0
0
7 Pulser~
4 153 395 0 10 12
0 72 73 74 46 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4460 0 0
2
5.89916e-315 0
0
5 4027~
219 356 434 0 7 32
0 75 15 46 15 76 11 12
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3260 0 0
2
5.89916e-315 5.42933e-315
0
5 4027~
219 488 432 0 7 32
0 18 13 11 13 77 10 16
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
5156 0 0
2
5.89916e-315 5.42414e-315
0
5 4027~
219 614 430 0 7 32
0 78 14 10 14 79 43 17
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U7A
12 -62 33 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
3133 0 0
2
5.89916e-315 5.41896e-315
0
79
7 7 3 0 0 4224 0 3 37 0 0 3
1137 467
1247 467
1247 434
8 6 4 0 0 4224 0 3 37 0 0 3
1137 476
1241 476
1241 434
9 5 5 0 0 4224 0 3 37 0 0 3
1137 485
1235 485
1235 434
10 4 6 0 0 4224 0 3 37 0 0 3
1137 494
1229 494
1229 434
11 3 7 0 0 4224 0 3 37 0 0 3
1137 503
1223 503
1223 434
12 2 8 0 0 4224 0 3 37 0 0 3
1137 512
1217 512
1217 434
1 13 9 0 0 4224 0 37 3 0 0 3
1211 434
1211 521
1137 521
0 3 10 0 0 4096 0 0 43 69 0 4
518 424
562 424
562 403
590 403
6 3 11 0 0 4096 0 41 42 0 0 4
386 416
425 416
425 405
464 405
0 7 12 0 0 4096 0 0 41 72 0 3
404 401
380 401
380 398
0 0 13 0 0 4224 0 0 0 17 75 4
472 714
472 449
459 449
459 414
0 0 14 0 0 4224 0 0 0 19 76 2
578 275
578 394
0 0 15 0 0 4224 0 0 0 0 79 3
308 505
308 416
316 416
0 4 12 0 0 8192 0 0 3 72 0 5
861 464
861 428
1018 428
1018 494
1073 494
0 3 16 0 0 8192 0 0 3 70 0 5
849 519
849 502
1064 502
1064 485
1073 485
0 2 17 0 0 8192 0 0 3 68 0 5
869 589
869 558
1045 558
1045 476
1073 476
5 0 13 0 0 128 0 32 0 0 0 2
477 714
468 714
0 1 18 0 0 8320 0 0 42 0 0 3
491 374
491 375
488 375
1 0 14 0 0 128 0 4 0 0 0 4
518 275
588 275
588 277
587 277
1 0 19 0 0 4224 0 5 0 0 0 3
258 507
324 506
324 504
1 3 20 0 0 8320 0 6 7 0 0 3
681 1099
681 1103
730 1103
1 3 21 0 0 8320 0 8 11 0 0 3
689 1199
689 1203
739 1203
3 1 22 0 0 8320 0 10 11 0 0 3
813 1240
790 1240
790 1212
3 2 23 0 0 4224 0 9 11 0 0 3
817 1172
790 1172
790 1194
1 3 24 0 0 8320 0 12 14 0 0 3
420 1090
420 1094
469 1094
3 2 25 0 0 8320 0 13 14 0 0 3
543 1061
520 1061
520 1085
1 0 12 0 0 0 0 17 0 0 72 3
737 341
778 341
778 464
2 0 26 0 0 4096 0 17 0 0 66 2
737 323
949 323
1 0 16 0 0 8192 0 15 0 0 70 3
736 279
824 279
824 519
2 0 26 0 0 4096 0 15 0 0 66 2
736 261
949 261
1 0 17 0 0 8320 0 16 0 0 68 3
732 225
791 225
791 589
2 0 27 0 0 4096 0 16 0 0 65 2
732 207
984 207
1 0 26 0 0 0 0 33 0 0 66 2
984 120
949 120
1 1 28 0 0 8320 0 3 1 0 0 4
1073 467
1053 467
1053 441
1052 441
1 2 29 0 0 4096 0 18 18 0 0 2
638 288
638 279
2 3 29 0 0 8320 0 18 17 0 0 4
638 279
680 279
680 332
686 332
3 3 30 0 0 4224 0 15 18 0 0 4
685 270
637 270
637 270
638 270
3 4 31 0 0 8320 0 16 18 0 0 4
681 216
637 216
637 261
638 261
1 3 32 0 0 8320 0 27 26 0 0 3
114 1118
114 1122
161 1122
3 1 33 0 0 4224 0 24 26 0 0 3
238 1164
238 1131
212 1131
3 2 34 0 0 4224 0 25 26 0 0 4
236 1091
211 1091
211 1113
212 1113
1 0 35 0 0 4096 0 22 0 0 43 3
215 997
225 997
225 988
2 3 35 0 0 8320 0 22 21 0 0 4
215 988
238 988
238 1043
249 1043
3 3 36 0 0 4224 0 22 20 0 0 4
215 979
242 979
242 994
248 994
4 3 37 0 0 4224 0 22 19 0 0 4
215 970
241 970
241 946
247 946
1 5 38 0 0 8320 0 23 22 0 0 3
116 980
116 984
164 984
0 2 17 0 0 0 0 0 28 51 0 3
691 697
691 765
633 765
0 1 12 0 0 0 0 0 28 49 0 3
657 740
657 783
633 783
0 1 12 0 0 4096 0 0 30 72 0 3
763 464
763 740
634 740
0 2 27 0 0 0 0 0 30 52 0 3
664 679
664 722
634 722
1 0 17 0 0 0 0 29 0 0 68 3
636 697
766 697
766 589
2 0 27 0 0 4096 0 29 0 0 65 2
636 679
985 679
1 0 11 0 0 8192 0 31 0 0 71 3
638 652
744 652
744 482
2 0 16 0 0 0 0 31 0 0 70 3
638 643
708 643
708 519
0 0 26 0 0 4096 0 0 0 60 66 2
638 629
949 629
5 4 39 0 0 8320 0 31 32 0 0 4
587 639
543 639
543 700
528 700
2 3 40 0 0 4224 0 32 30 0 0 4
528 718
577 718
577 731
583 731
3 3 41 0 0 4224 0 29 32 0 0 4
585 688
538 688
538 709
528 709
3 1 42 0 0 8320 0 28 32 0 0 4
582 774
538 774
538 727
528 727
4 3 26 0 0 0 0 31 31 0 0 2
638 625
638 634
6 0 43 0 0 12416 0 43 0 0 0 4
644 412
643 412
643 612
877 612
1 0 43 0 0 0 0 35 0 0 61 2
457 545
643 545
2 0 27 0 0 0 0 35 0 0 64 2
457 527
457 495
2 0 27 0 0 4224 0 34 0 0 65 2
375 495
985 495
2 0 27 0 0 0 0 33 0 0 0 4
984 156
984 495
985 495
985 913
1 0 26 0 0 4224 0 2 0 0 0 2
949 107
949 913
3 1 44 0 0 8320 0 35 34 0 0 4
406 536
388 536
388 513
375 513
7 0 17 0 0 0 0 43 0 0 0 4
638 394
662 394
662 589
877 589
6 0 10 0 0 8320 0 42 0 0 0 3
518 414
518 539
873 539
7 0 16 0 0 12416 0 42 0 0 0 4
512 396
522 396
522 519
873 519
6 0 11 0 0 8320 0 41 0 0 0 3
386 416
386 482
875 482
0 0 12 0 0 8320 0 0 0 0 0 3
404 398
404 464
877 464
1 9 2 0 0 4224 0 36 37 0 0 2
1232 335
1232 356
1 3 45 0 0 8320 0 38 0 0 0 3
91 233
91 237
138 237
2 4 13 0 0 128 0 42 42 0 0 4
464 396
454 396
454 414
464 414
2 4 14 0 0 128 0 43 43 0 0 4
590 394
578 394
578 412
590 412
1 0 46 0 0 4096 0 39 0 0 78 2
193 329
193 407
3 4 46 0 0 4224 0 41 40 0 0 3
332 407
183 407
183 395
2 4 15 0 0 128 0 41 41 0 0 4
332 398
313 398
313 416
332 416
17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
625 342 654 366
635 350 643 366
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
505 344 534 368
515 352 523 368
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
875 444 904 468
885 452 893 468
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
872 465 909 489
882 473 898 489
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
870 500 899 524
880 508 888 524
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
872 522 909 546
882 530 898 546
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
874 569 903 593
884 577 892 593
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
875 593 912 617
885 601 901 617
2 C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
295 476 332 500
305 484 321 500
2 Ta
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
462 684 499 708
472 692 488 708
2 Tb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
147 1092 184 1116
157 1100 173 1116
2 Kb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
148 955 185 979
158 963 174 979
2 Jb
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
424 1054 485 1078
434 1062 474 1078
5 Ja,Ka
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
719 1173 756 1197
729 1181 745 1197
2 Jc
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
719 1073 756 1097
729 1081 745 1097
2 Kc
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
567 247 604 271
577 255 593 271
2 Tc
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
375 349 404 373
385 357 393 373
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
