CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 147 243 0 1 11
0 17
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
5.89912e-315 5.32571e-315
0
13 Logic Switch~
5 119 242 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3820 0 0
2
5.89912e-315 5.30499e-315
0
13 Logic Switch~
5 89 242 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
5.89912e-315 5.26354e-315
0
13 Logic Switch~
5 55 241 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
5.89912e-315 0
0
5 SCOPE
12 450 156 0 1 11
0 3
0
0 0 57584 0
3 TP7
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3178 0 0
2
5.89912e-315 0
0
5 SCOPE
12 770 235 0 1 11
0 4
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3409 0 0
2
5.89912e-315 0
0
5 SCOPE
12 503 232 0 1 11
0 3
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3951 0 0
2
5.89912e-315 0
0
5 SCOPE
12 639 233 0 1 11
0 5
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8885 0 0
2
5.89912e-315 0
0
5 SCOPE
12 1025 587 0 1 11
0 6
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3780 0 0
2
5.89912e-315 0
0
5 SCOPE
12 949 308 0 1 11
0 7
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9265 0 0
2
5.89912e-315 0
0
5 SCOPE
12 352 256 0 1 11
0 8
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9442 0 0
2
5.89912e-315 0
0
14 Logic Display~
6 1061 485 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89912e-315 0
0
14 Logic Display~
6 587 436 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.89912e-315 5.26354e-315
0
14 Logic Display~
6 441 437 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89912e-315 0
0
14 Logic Display~
6 712 437 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89912e-315 5.26354e-315
0
14 Logic Display~
6 816 436 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89912e-315 0
0
6 74LS85
106 923 562 0 14 29
0 14 15 16 17 12 10 11 9 20
21 22 23 13 6
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U1
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3171 0 0
2
5.89912e-315 0
0
9 Inverter~
13 1001 337 0 2 22
0 13 7
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U4A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4139 0 0
2
5.89912e-315 0
0
2 +V
167 344 85 0 1 3
0 19
0
0 0 54256 0
2 5V
-7 -21 7 -13
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
5.89912e-315 0
0
7 Pulser~
4 312 277 0 10 12
0 2 2 8 24 0 0 5 5 4
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5283 0 0
2
5.89912e-315 5.43192e-315
0
5 7474~
219 831 269 0 6 22
0 19 18 4 7 18 12
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U3B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 2 0
1 U
6874 0 0
2
5.89912e-315 5.42933e-315
0
5 7474~
219 698 265 0 6 22
0 19 4 5 7 4 10
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 2 0
1 U
5305 0 0
2
5.89912e-315 5.42414e-315
0
5 7474~
219 564 263 0 6 22
0 19 5 3 7 5 11
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 1 0
1 U
34 0 0
2
5.89912e-315 5.41896e-315
0
5 7474~
219 424 262 0 6 22
0 19 3 8 7 3 9
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 1 0
1 U
969 0 0
2
5.89912e-315 5.41378e-315
0
7 Ground~
168 220 287 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8402 0 0
2
5.89912e-315 5.4086e-315
0
39
1 0 3 0 0 0 0 5 0 0 33 2
450 168
450 168
1 0 4 0 0 0 0 6 0 0 34 2
770 247
770 247
1 0 3 0 0 0 0 7 0 0 36 2
503 244
503 244
1 0 5 0 0 0 0 8 0 0 35 2
639 245
639 245
1 0 6 0 0 4096 0 9 0 0 8 2
1025 599
1025 598
1 0 7 0 0 4096 0 10 0 0 28 2
949 320
949 319
1 0 8 0 0 0 0 11 0 0 37 2
352 268
352 268
14 1 6 0 0 4224 0 17 12 0 0 3
955 598
1061 598
1061 503
6 0 9 0 0 8192 0 24 0 0 13 3
448 226
463 226
463 509
6 0 10 0 0 8192 0 22 0 0 16 3
722 229
741 229
741 486
6 0 11 0 0 8192 0 23 0 0 15 3
588 227
604 227
604 499
6 0 12 0 0 8192 0 21 0 0 17 3
855 233
865 233
865 472
8 1 9 0 0 20608 0 17 14 0 0 7
891 598
679 598
679 651
959 651
959 509
441 509
441 455
13 1 13 0 0 8320 0 17 18 0 0 5
955 589
1097 589
1097 381
1004 381
1004 355
7 1 11 0 0 20608 0 17 13 0 0 7
891 589
660 589
660 665
971 665
971 499
587 499
587 454
6 1 10 0 0 12416 0 17 15 0 0 7
891 580
640 580
640 686
989 686
989 486
712 486
712 455
5 1 12 0 0 12416 0 17 16 0 0 7
891 571
624 571
624 700
1005 700
1005 472
816 472
816 454
1 1 14 0 0 4224 0 17 4 0 0 3
891 535
55 535
55 253
2 1 15 0 0 4224 0 17 3 0 0 3
891 544
89 544
89 254
3 1 16 0 0 4224 0 17 2 0 0 3
891 553
119 553
119 254
4 1 17 0 0 4224 0 17 1 0 0 3
891 562
147 562
147 255
2 5 18 0 0 12416 0 21 21 0 0 6
807 233
790 233
790 175
883 175
883 251
861 251
2 0 4 0 0 12416 0 22 0 0 34 5
674 229
662 229
662 189
751 189
751 247
2 0 5 0 0 12416 0 23 0 0 35 5
540 227
531 227
531 189
614 189
614 245
4 0 7 0 0 4096 0 21 0 0 28 2
831 281
831 319
4 0 7 0 0 4096 0 22 0 0 28 2
698 277
698 319
4 0 7 0 0 4096 0 23 0 0 28 2
564 275
564 319
2 4 7 0 0 4224 0 18 24 0 0 3
1004 319
424 319
424 274
1 0 19 0 0 4096 0 22 0 0 32 2
698 202
698 134
1 0 19 0 0 0 0 23 0 0 32 2
564 200
564 134
1 0 19 0 0 0 0 24 0 0 32 2
424 199
424 134
1 1 19 0 0 8320 0 19 21 0 0 4
344 94
344 134
831 134
831 206
2 0 3 0 0 12416 0 24 0 0 36 5
400 226
378 226
378 168
477 168
477 244
5 3 4 0 0 0 0 22 21 0 0 4
728 247
799 247
799 251
807 251
5 3 5 0 0 0 0 23 22 0 0 4
594 245
666 245
666 247
674 247
5 3 3 0 0 0 0 24 23 0 0 4
454 244
532 244
532 245
540 245
3 3 8 0 0 4224 0 20 24 0 0 4
336 268
377 268
377 244
400 244
2 0 2 0 0 4096 0 20 0 0 39 3
282 277
255 277
255 268
1 1 2 0 0 4224 0 20 25 0 0 3
288 268
220 268
220 281
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
64 35 157 59
74 43 146 59
9 Quest�o 2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
