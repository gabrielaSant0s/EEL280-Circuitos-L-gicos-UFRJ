CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 70 1 90 10
172 80 1364 539
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 2 0.253589 0.500000
172 548 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 667 445 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 180
2 5V
16 1 30 9
2 Q2
17 -11 31 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.89912e-315 0
0
13 Logic Switch~
5 668 408 0 1 11
0 11
0
0 0 21360 180
2 0V
16 3 30 11
2 Q3
15 -7 29 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
5.89912e-315 0
0
13 Logic Switch~
5 665 523 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 180
2 5V
16 2 30 10
2 Q0
15 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
5.89912e-315 5.32571e-315
0
13 Logic Switch~
5 666 485 0 1 11
0 9
0
0 0 21360 180
2 0V
15 4 29 12
2 Q1
15 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
5.89912e-315 5.30499e-315
0
13 Logic Switch~
5 399 118 0 1 11
0 25
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 UD
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
5.89912e-315 0
0
13 Logic Switch~
5 430 119 0 1 11
0 26
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 CE
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3178 0 0
2
5.89912e-315 0
0
5 SCOPE
12 720 202 0 1 11
0 3
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3409 0 0
2
43759.4 0
0
5 SCOPE
12 695 220 0 1 11
0 4
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3951 0 0
2
43759.4 0
0
5 SCOPE
12 666 236 0 1 11
0 5
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8885 0 0
2
43759.4 0
0
5 SCOPE
12 635 257 0 1 11
0 6
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3780 0 0
2
43759.4 0
0
5 SCOPE
12 419 317 0 1 11
0 2
0
0 0 57584 90
3 TP2
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9265 0 0
2
43759.4 1
0
5 SCOPE
12 302 244 0 1 11
0 7
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9442 0 0
2
43759.4 0
0
10 2-In XNOR~
219 509 514 0 3 22
0 8 3 12
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4D
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
9424 0 0
2
5.89912e-315 0
0
10 2-In XNOR~
219 510 477 0 3 22
0 9 4 13
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4C
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
9968 0 0
2
5.89912e-315 0
0
10 2-In XNOR~
219 511 436 0 3 22
0 10 5 14
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4B
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9281 0 0
2
5.89912e-315 0
0
10 2-In XNOR~
219 511 399 0 3 22
0 11 6 15
0
0 0 624 180
4 4077
-7 -24 21 -16
3 U4A
4 -25 25 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
8464 0 0
2
5.89912e-315 0
0
5 7422~
219 429 446 0 5 22
0 12 14 13 15 16
0
0 0 624 180
6 74LS22
-21 -28 21 -20
3 U3A
-8 -31 13 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
7168 0 0
2
5.89912e-315 0
0
2 +V
167 834 151 0 1 3
0 17
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3171 0 0
2
5.89912e-315 0
0
9 CA 7-Seg~
184 834 194 0 18 19
10 24 23 22 21 20 19 18 27 17
0 0 2 0 0 2 0 2 1
0
0 0 21088 0
8 YELLOWCA
6 -41 62 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4139 0 0
2
5.89912e-315 0
0
7 Ground~
168 429 337 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
5.89912e-315 0
0
14 Logic Display~
6 235 193 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.89912e-315 0
0
7 Pulser~
4 160 264 0 10 12
0 28 29 7 30 0 0 5 5 4
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6874 0 0
2
5.89912e-315 0
0
6 74LS47
187 763 319 0 14 29
0 6 5 4 3 31 32 18 19 20
21 22 23 24 33
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5305 0 0
2
5.89912e-315 0
0
7 74LS190
134 480 273 0 14 29
0 26 7 16 25 2 2 2 2 34
35 6 5 4 3
0
0 0 4848 0
6 74F190
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
5.89912e-315 0
0
40
1 0 3 0 0 4096 0 7 0 0 35 2
720 214
720 310
1 0 4 0 0 4096 0 8 0 0 36 2
695 232
695 301
1 0 5 0 0 4096 0 9 0 0 37 2
666 248
666 292
1 0 6 0 0 4096 0 10 0 0 38 2
635 269
635 283
1 0 2 0 0 0 0 11 0 0 34 2
429 319
429 319
8 0 2 0 0 4096 0 24 0 0 34 2
448 309
429 309
1 0 7 0 0 4096 0 12 0 0 39 2
302 256
302 255
1 1 8 0 0 4224 0 13 3 0 0 2
537 523
651 523
1 1 9 0 0 4224 0 14 4 0 0 3
538 486
652 486
652 485
1 1 10 0 0 4224 0 15 1 0 0 2
539 445
653 445
1 1 11 0 0 4224 0 16 2 0 0 2
539 408
654 408
2 0 3 0 0 8320 0 13 0 0 35 3
537 505
631 505
631 309
2 0 4 0 0 8320 0 14 0 0 36 3
538 468
603 468
603 300
2 0 5 0 0 8192 0 15 0 0 37 3
539 427
578 427
578 291
2 0 6 0 0 8192 0 16 0 0 38 3
539 390
553 390
553 282
1 3 12 0 0 8320 0 17 13 0 0 4
453 464
468 464
468 514
482 514
3 3 13 0 0 4224 0 17 14 0 0 3
453 452
483 452
483 477
2 3 14 0 0 4224 0 17 15 0 0 3
453 440
484 440
484 436
4 3 15 0 0 8320 0 17 16 0 0 4
453 428
464 428
464 399
484 399
3 5 16 0 0 8320 0 24 17 0 0 4
442 264
349 264
349 446
402 446
1 9 17 0 0 4224 0 18 19 0 0 2
834 160
834 158
7 7 18 0 0 8320 0 23 19 0 0 3
801 283
849 283
849 230
8 6 19 0 0 8320 0 23 19 0 0 3
801 292
843 292
843 230
9 5 20 0 0 8320 0 23 19 0 0 3
801 301
837 301
837 230
10 4 21 0 0 8320 0 23 19 0 0 3
801 310
831 310
831 230
11 3 22 0 0 8320 0 23 19 0 0 3
801 319
825 319
825 230
12 2 23 0 0 8320 0 23 19 0 0 3
801 328
819 328
819 230
13 1 24 0 0 8320 0 23 19 0 0 3
801 337
813 337
813 230
1 0 25 0 0 0 0 5 0 0 30 2
399 130
399 130
4 0 25 0 0 8320 0 24 0 0 0 3
448 273
399 273
399 127
1 1 26 0 0 4224 0 6 24 0 0 3
430 131
430 246
442 246
7 0 2 0 0 0 0 24 0 0 34 2
448 300
429 300
6 0 2 0 0 0 0 24 0 0 34 2
448 291
429 291
1 5 2 0 0 4224 0 20 24 0 0 3
429 331
429 282
448 282
14 4 3 0 0 0 0 24 23 0 0 4
512 309
631 309
631 310
731 310
13 3 4 0 0 0 0 24 23 0 0 4
512 300
603 300
603 301
731 301
12 2 5 0 0 12416 0 24 23 0 0 4
512 291
578 291
578 292
731 292
11 1 6 0 0 12416 0 24 23 0 0 4
512 282
553 282
553 283
731 283
0 2 7 0 0 4224 0 0 24 40 0 2
235 255
448 255
3 1 7 0 0 0 0 22 21 0 0 3
184 255
235 255
235 211
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
