CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 550 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
61
2 +V
167 305 1155 0 1 3
0 0
0
0 0 54240 0
2 5V
-8 -22 6 -14
3 VCC
-9 -34 12 -26
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3805 0 0
2
43739.1 0
0
13 Logic Switch~
5 109 1684 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 D
-20 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5219 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 109 1658 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 C
-21 -5 -14 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3795 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 109 1630 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 B
-20 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3637 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 109 1600 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 A
-20 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3226 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 68 1384 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
29 -12 43 -4
1 D
12 -11 19 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6966 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 66 1345 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
36 -11 50 -3
1 C
19 -10 26 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9796 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 69 1317 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
16 -11 30 -3
1 B
-2 -15 5 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5952 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 79 1283 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
32 -13 46 -5
1 A
19 -13 26 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3649 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 334 1418 0 1 11
0 30
0
0 0 21344 0
2 0V
9 4 23 12
2 V3
10 -10 24 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3716 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 335 1400 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
12 -12 26 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4797 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 271 629 0 1 11
0 43
0
0 0 21344 270
2 0V
-7 -20 7 -12
2 D1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4681 0 0
2
43739.1 0
0
13 Logic Switch~
5 102 631 0 1 11
0 41
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9730 0 0
2
43739.1 1
0
13 Logic Switch~
5 150 631 0 1 11
0 38
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9874 0 0
2
43739.1 2
0
13 Logic Switch~
5 208 629 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-7 -20 7 -12
2 C1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
364 0 0
2
43739.1 3
0
13 Logic Switch~
5 214 87 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3656 0 0
2
5.8991e-315 0
0
13 Logic Switch~
5 157 88 0 10 11
0 54 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3131 0 0
2
5.8991e-315 5.26354e-315
0
13 Logic Switch~
5 105 90 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6772 0 0
2
5.8991e-315 5.30499e-315
0
5 4023~
219 752 1951 0 4 22
0 4 6 5 3
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U16B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 16 0
1 U
9557 0 0
2
5.8991e-315 0
0
5 4012~
219 662 1993 0 5 22
0 10 9 8 7 5
0
0 0 608 0
4 4012
-7 -24 21 -16
4 U17A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 17 0
1 U
5789 0 0
2
5.8991e-315 0
0
5 4012~
219 563 1937 0 5 22
0 10 12 11 7 6
0
0 0 608 0
4 4012
-7 -24 21 -16
4 U15B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 2 15 0
1 U
7328 0 0
2
5.8991e-315 0
0
5 4023~
219 435 1886 0 4 22
0 4 15 14 13
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U16A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 16 0
1 U
4799 0 0
2
5.8991e-315 0
0
5 4012~
219 333 1912 0 5 22
0 16 11 9 17 14
0
0 0 608 0
4 4012
-7 -24 21 -16
4 U15A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 15 0
1 U
9196 0 0
2
5.8991e-315 0
0
5 4012~
219 333 1863 0 5 22
0 16 8 9 17 15
0
0 0 608 0
4 4012
-7 -24 21 -16
4 U14B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 2 14 0
1 U
3857 0 0
2
5.8991e-315 0
0
5 4012~
219 234 1812 0 5 22
0 7 11 9 17 4
0
0 0 608 0
4 4012
-7 -24 21 -16
4 U14A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 14 0
1 U
7125 0 0
2
5.8991e-315 0
0
5 4049~
219 224 1767 0 2 22
0 7 16
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U12E
6 -13 34 -5
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 11 0
1 U
3641 0 0
2
5.8991e-315 0
0
5 4049~
219 224 1748 0 2 22
0 11 8
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U12D
10 -12 38 -4
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 11 0
1 U
9821 0 0
2
5.8991e-315 0
0
5 4049~
219 224 1729 0 2 22
0 9 12
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U12C
5 -14 33 -6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 11 0
1 U
3187 0 0
2
5.8991e-315 0
0
5 4049~
219 223 1709 0 2 22
0 17 10
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U12B
6 -14 34 -6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
762 0 0
2
5.8991e-315 0
0
14 Logic Display~
6 851 1611 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
39 0 0
2
5.8991e-315 0
0
14 Logic Display~
6 825 1611 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9450 0 0
2
5.8991e-315 0
0
14 Logic Display~
6 792 1612 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3236 0 0
2
5.8991e-315 0
0
14 Logic Display~
6 611 1300 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3321 0 0
2
5.8991e-315 0
0
14 Logic Display~
6 677 1302 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8879 0 0
2
5.8991e-315 0
0
14 Logic Display~
6 753 1304 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5433 0 0
2
5.8991e-315 0
0
8 3-In OR~
219 476 1444 0 4 22
0 21 20 19 18
0
0 0 608 0
4 4075
-14 -24 14 -16
4 U13B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 13 0
1 U
3679 0 0
2
5.8991e-315 0
0
8 3-In OR~
219 466 1371 0 4 22
0 21 24 23 22
0
0 0 608 0
4 4075
-14 -24 14 -16
4 U13A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 13 0
1 U
9342 0 0
2
5.8991e-315 0
0
5 4049~
219 466 1328 0 2 22
0 21 25
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U12A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
3623 0 0
2
5.8991e-315 0
0
4 4514
219 393 1391 0 30 45
0 29 28 27 26 31 30 56 57 58
19 59 20 60 61 62 63 64 65 23
66 24 21 0 0 0 0 0 0 0
15
0
0 0 4832 0
4 4514
-14 -87 14 -79
3 U10
-11 -88 10 -80
0
16 DVDD=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 22 21 3 2 1 23 11 9 10
8 7 6 5 4 18 17 20 19 14
13 16 15 22 21 3 2 1 23 11
9 10 8 7 6 5 4 18 17 20
19 14 13 16 15 0
65 0 0 512 1 0 0 0
1 U
3722 0 0
2
5.8991e-315 0
0
5 4023~
219 527 1035 0 4 22
0 36 35 34 33
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U11C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 12 0
1 U
8993 0 0
2
43739.1 4
0
5 4023~
219 322 1073 0 4 22
0 32 32 67 37
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U11B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 512 3 2 12 0
1 U
3723 0 0
2
43739.1 5
0
5 4023~
219 411 1094 0 4 22
0 39 38 37 34
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U11A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 12 0
1 U
6244 0 0
2
43739.1 6
0
10 2-In NAND~
219 410 1035 0 3 22
0 40 32 35
0
0 0 608 0
6 74LS37
-14 -24 28 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
6421 0 0
2
43739.1 7
0
10 2-In NAND~
219 412 980 0 3 22
0 41 40 36
0
0 0 608 0
6 74LS37
-14 -24 28 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
7743 0 0
2
43739.1 8
0
14 Logic Display~
6 603 1015 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9840 0 0
2
43739.1 9
0
10 2-In NAND~
219 319 1007 0 3 22
0 38 38 40
0
0 0 608 0
6 74LS37
-14 -24 28 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
6910 0 0
2
43739.1 10
0
10 2-In NAND~
219 323 945 0 3 22
0 41 41 39
0
0 0 608 0
6 74LS37
-14 -24 28 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
449 0 0
2
43739.1 11
0
14 Logic Display~
6 693 732 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8761 0 0
2
43739.1 12
0
7 Ground~
168 602 711 0 1 3
0 2
0
0 0 53344 692
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6748 0 0
2
43739.1 13
0
7 74LS153
119 507 772 0 14 29
0 44 45 44 45 38 43 68 69 70
71 2 72 42 73
0
0 0 4832 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
7393 0 0
2
43739.1 14
0
9 Inverter~
13 400 762 0 2 22
0 44 45
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
7699 0 0
2
43739.1 15
0
5 7433~
219 317 720 0 3 22
0 41 32 44
0
0 0 608 0
6 74LS33
-21 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 2 3 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6638 0 0
2
43739.1 16
0
14 Logic Display~
6 439 484 0 1 2
10 48
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
5.8991e-315 5.32571e-315
0
10 2-In NAND~
219 376 506 0 3 22
0 47 46 48
0
0 0 608 0
5 74F37
-10 -24 25 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
9395 0 0
2
5.8991e-315 5.34643e-315
0
14 Logic Display~
6 656 297 0 1 2
10 49
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3303 0 0
2
5.8991e-315 5.3568e-315
0
10 2-In NAND~
219 600 315 0 3 22
0 51 50 49
0
0 0 608 0
5 74F37
-10 -24 25 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
4498 0 0
2
5.8991e-315 5.36716e-315
0
5 7433~
219 507 393 0 3 22
0 53 52 50
0
0 0 608 0
6 74LS33
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 2 3 1 2 3 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9728 0 0
2
5.8991e-315 5.37752e-315
0
8 2-In OR~
219 490 242 0 3 22
0 47 53 51
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3789 0 0
2
5.8991e-315 5.38788e-315
0
9 3-In NOR~
219 423 323 0 4 22
0 52 54 47 53
0
0 0 608 0
5 74F27
-18 -24 17 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
3978 0 0
2
5.8991e-315 5.39306e-315
0
9 2-In XOR~
219 328 284 0 3 22
0 46 55 52
0
0 0 608 0
5 74F86
-18 -24 17 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3494 0 0
2
5.8991e-315 5.39824e-315
0
2 +V
167 271 79 0 1 3
0 55
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3507 0 0
2
5.8991e-315 5.40342e-315
0
110
2 0 0 0 0 0 0 43 0 0 7 2
386 1044
365 1044
1 0 0 0 0 0 0 43 0 0 89 2
386 1026
208 1026
3 0 0 0 0 0 0 42 0 0 88 2
387 1103
271 1103
3 2 0 0 0 0 0 46 42 0 0 4
346 1007
353 1007
353 1094
387 1094
3 1 0 0 0 0 0 47 42 0 0 4
350 945
377 945
377 1085
387 1085
1 0 0 0 0 0 0 44 0 0 91 2
388 971
102 971
4 2 0 0 0 0 0 41 44 0 0 4
349 1073
365 1073
365 989
388 989
2 0 0 0 0 0 0 41 0 0 9 3
298 1073
286 1073
286 1064
1 0 0 0 0 0 0 41 0 0 88 2
298 1064
271 1064
2 0 0 0 0 0 0 46 0 0 11 3
295 1016
286 1016
286 998
1 0 0 0 0 0 0 46 0 0 89 2
295 998
208 998
3 1 0 0 0 0 0 41 1 0 0 5
298 1082
288 1082
288 1183
305 1183
305 1164
4 1 3 0 0 8320 0 19 32 0 0 3
779 1951
792 1951
792 1630
1 0 4 0 0 8192 0 19 0 0 37 3
728 1942
722 1942
722 1812
3 5 5 0 0 8320 0 19 20 0 0 4
728 1960
705 1960
705 1993
689 1993
5 2 6 0 0 4224 0 21 19 0 0 4
590 1937
704 1937
704 1951
728 1951
4 0 7 0 0 8192 0 20 0 0 50 3
638 2007
604 2007
604 1684
3 0 8 0 0 8192 0 20 0 0 43 3
638 1998
615 1998
615 1748
2 0 9 0 0 8192 0 20 0 0 52 3
638 1989
632 1989
632 1630
1 0 10 0 0 8192 0 20 0 0 45 3
638 1980
623 1980
623 1709
4 0 7 0 0 0 0 21 0 0 50 3
539 1951
518 1951
518 1684
3 0 11 0 0 8192 0 21 0 0 51 3
539 1942
503 1942
503 1658
2 0 12 0 0 8192 0 21 0 0 44 3
539 1933
481 1933
481 1729
0 1 10 0 0 0 0 0 21 45 0 3
489 1709
489 1924
539 1924
4 1 13 0 0 4224 0 22 31 0 0 3
462 1886
825 1886
825 1629
1 0 4 0 0 0 0 22 0 0 37 3
411 1877
387 1877
387 1812
5 3 14 0 0 12416 0 23 22 0 0 4
360 1912
379 1912
379 1895
411 1895
5 2 15 0 0 12416 0 24 22 0 0 4
360 1863
378 1863
378 1886
411 1886
0 1 16 0 0 4096 0 0 23 33 0 3
283 1850
283 1899
309 1899
2 0 11 0 0 0 0 23 0 0 40 3
309 1908
183 1908
183 1808
3 0 9 0 0 0 0 23 0 0 35 3
309 1917
158 1917
158 1868
0 4 17 0 0 8192 0 0 23 36 0 3
134 1877
134 1926
309 1926
1 0 16 0 0 8192 0 24 0 0 42 3
309 1850
269 1850
269 1767
0 2 8 0 0 0 0 0 24 43 0 3
261 1748
261 1859
309 1859
3 0 9 0 0 0 0 24 0 0 39 3
309 1868
158 1868
158 1817
0 4 17 0 0 0 0 0 24 38 0 3
134 1826
134 1877
309 1877
5 1 4 0 0 4224 0 25 30 0 0 3
261 1812
851 1812
851 1629
0 4 17 0 0 0 0 0 25 49 0 3
134 1709
134 1826
210 1826
3 0 9 0 0 0 0 25 0 0 48 3
210 1817
158 1817
158 1729
2 0 11 0 0 0 0 25 0 0 47 3
210 1808
182 1808
182 1748
0 1 7 0 0 0 0 0 25 46 0 3
199 1765
199 1799
210 1799
2 0 16 0 0 4224 0 26 0 0 0 2
245 1767
707 1767
2 0 8 0 0 4224 0 27 0 0 0 2
245 1748
707 1748
2 0 12 0 0 4224 0 28 0 0 0 2
245 1729
707 1729
2 0 10 0 0 4224 0 29 0 0 0 2
244 1709
707 1709
0 1 7 0 0 0 0 0 26 50 0 3
199 1684
199 1767
209 1767
0 1 11 0 0 0 0 0 27 51 0 3
182 1658
182 1748
209 1748
0 1 9 0 0 0 0 0 28 52 0 3
158 1630
158 1729
209 1729
0 1 17 0 0 0 0 0 29 53 0 3
134 1600
134 1709
208 1709
1 0 7 0 0 4224 0 2 0 0 0 2
121 1684
707 1684
1 0 11 0 0 4224 0 3 0 0 0 2
121 1658
706 1658
1 0 9 0 0 4224 0 4 0 0 0 2
121 1630
707 1630
1 0 17 0 0 4224 0 5 0 0 0 2
121 1600
709 1600
4 1 18 0 0 8320 0 36 33 0 0 3
509 1444
611 1444
611 1318
10 3 19 0 0 12416 0 39 36 0 0 4
425 1436
435 1436
435 1453
463 1453
2 12 20 0 0 8320 0 36 39 0 0 4
464 1444
442 1444
442 1418
425 1418
0 1 21 0 0 4224 0 0 36 61 0 3
448 1362
448 1435
463 1435
4 1 22 0 0 4224 0 37 34 0 0 3
499 1371
677 1371
677 1320
19 3 23 0 0 8320 0 39 37 0 0 4
425 1355
436 1355
436 1380
453 1380
2 21 24 0 0 8320 0 37 39 0 0 4
454 1371
442 1371
442 1337
425 1337
1 0 21 0 0 0 0 37 0 0 63 3
453 1362
447 1362
447 1328
2 1 25 0 0 4224 0 38 35 0 0 3
487 1328
753 1328
753 1322
22 1 21 0 0 0 0 39 38 0 0 2
425 1328
451 1328
1 4 26 0 0 4224 0 6 39 0 0 4
80 1384
269 1384
269 1373
361 1373
1 3 27 0 0 4224 0 7 39 0 0 4
78 1345
290 1345
290 1364
361 1364
1 2 28 0 0 12416 0 8 39 0 0 6
81 1317
82 1317
82 1318
302 1318
302 1355
361 1355
1 1 29 0 0 4224 0 9 39 0 0 4
91 1283
313 1283
313 1346
361 1346
1 6 30 0 0 12416 0 10 39 0 0 4
346 1418
343 1418
343 1418
355 1418
5 1 31 0 0 4224 0 39 11 0 0 2
361 1400
347 1400
4 1 33 0 0 4224 0 40 45 0 0 5
554 1035
591 1035
591 1041
603 1041
603 1033
4 3 34 0 0 8320 0 42 40 0 0 4
438 1094
455 1094
455 1044
503 1044
3 2 35 0 0 4224 0 43 40 0 0 2
437 1035
503 1035
3 1 36 0 0 12432 0 44 40 0 0 4
439 980
453 980
453 1026
503 1026
2 0 41 0 0 0 0 47 0 0 75 3
299 954
287 954
287 936
1 0 41 0 0 0 0 47 0 0 91 2
299 936
102 936
3 1 42 0 0 4096 0 0 48 77 0 3
657 754
693 754
693 750
13 0 42 0 0 4224 0 50 0 0 76 2
539 754
659 754
11 1 2 0 0 4224 0 50 49 0 0 3
545 736
602 736
602 719
6 0 43 0 0 4096 0 50 0 0 88 2
475 781
271 781
5 0 38 0 0 4096 0 50 0 0 90 2
475 772
150 772
3 0 44 0 0 4096 0 50 0 0 82 3
475 754
443 754
443 736
1 0 44 0 0 4224 0 50 0 0 85 2
475 736
372 736
2 0 45 0 0 4096 0 50 0 0 84 3
475 745
455 745
455 763
2 4 45 0 0 8320 0 51 50 0 0 3
421 762
421 763
475 763
3 1 44 0 0 0 0 52 51 0 0 4
356 720
372 720
372 762
385 762
2 0 32 0 0 0 0 52 0 0 89 2
304 729
208 729
1 0 41 0 0 0 0 52 0 0 91 2
304 711
102 711
1 0 43 0 0 4224 0 12 0 0 0 2
271 641
271 1179
1 0 32 0 0 4224 0 15 0 0 0 2
208 641
208 1179
1 0 38 0 0 4224 0 14 0 0 0 2
150 643
150 1180
1 0 41 0 0 4224 0 13 0 0 0 2
102 643
102 1179
2 0 46 0 0 4096 0 54 0 0 108 2
352 515
214 515
1 0 47 0 0 4096 0 54 0 0 110 2
352 497
105 497
3 1 48 0 0 4224 0 54 53 0 0 3
403 506
439 506
439 502
3 1 49 0 0 4224 0 56 55 0 0 2
627 315
656 315
3 2 50 0 0 8320 0 57 56 0 0 4
546 393
571 393
571 324
576 324
3 1 51 0 0 8320 0 58 56 0 0 4
523 242
571 242
571 306
576 306
0 2 52 0 0 8320 0 0 57 104 0 3
367 284
367 402
494 402
0 1 53 0 0 4096 0 0 57 101 0 3
469 323
469 384
494 384
1 0 47 0 0 4096 0 58 0 0 110 2
477 233
105 233
4 2 53 0 0 8320 0 59 58 0 0 4
462 323
469 323
469 251
477 251
3 0 47 0 0 0 0 59 0 0 110 2
410 332
105 332
2 0 54 0 0 4096 0 59 0 0 109 2
411 323
157 323
3 1 52 0 0 0 0 60 59 0 0 4
361 284
402 284
402 314
410 314
2 0 55 0 0 4096 0 60 0 0 107 2
312 293
271 293
1 0 46 0 0 0 0 60 0 0 108 2
312 275
214 275
1 0 55 0 0 4224 0 61 0 0 0 2
271 88
271 544
1 0 46 0 0 4224 0 16 0 0 0 2
214 99
214 545
1 0 54 0 0 4224 0 17 0 0 0 2
157 100
157 547
1 0 47 0 0 4224 0 18 0 0 0 2
105 102
105 547
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
345 431 582 455
355 439 571 455
27 LETRA A - CIRCUITO REDUZIDO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
362 169 599 193
372 177 588 193
27 LETRA A - CIRCUITO ORIGINAL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 28
386 892 631 916
396 900 620 916
28 LETRA B - CIRCUITO OTIMIZADO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
371 635 608 659
381 643 597 659
27 LETRA B - CIRCUITO ORIGINAL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
363 1232 528 1256
373 1240 517 1256
18 LETRA C - ORIGINAL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
369 1520 542 1544
379 1528 531 1544
19 LETRA C - OTIMIZADA
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
