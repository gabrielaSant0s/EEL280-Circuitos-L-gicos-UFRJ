CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 122 298 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43759 3
0
13 Logic Switch~
5 121 328 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43759 2
0
13 Logic Switch~
5 123 361 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43759 1
0
13 Logic Switch~
5 120 265 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43759 0
0
13 Logic Switch~
5 122 235 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43759 1
0
13 Logic Switch~
5 120 202 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43759 0
0
13 Logic Switch~
5 121 172 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43759 0
0
13 Logic Switch~
5 119 139 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43759 0
0
5 4049~
219 264 255 0 2 22
0 13 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
4747 0 0
2
43759 1
0
5 4049~
219 263 281 0 2 22
0 14 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
972 0 0
2
43759 0
0
5 4049~
219 264 230 0 2 22
0 12 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
3472 0 0
2
43759 0
0
5 4049~
219 265 204 0 2 22
0 11 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
9998 0 0
2
43759 0
0
7 Ground~
168 682 244 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
3536 0 0
2
43759 0
0
7 Ground~
168 323 58 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4597 0 0
2
43759 0
0
7 Ground~
168 595 81 0 1 3
0 2
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
3835 0 0
2
43759 0
0
7 Ground~
168 591 325 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3670 0 0
2
43759 0
0
8 3-In OR~
219 529 293 0 4 22
0 24 23 22 26
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 1 2 0
1 U
5616 0 0
2
43759 0
0
5 4081~
219 454 318 0 3 22
0 20 19 22
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9323 0 0
2
43759 0
0
5 4081~
219 452 264 0 3 22
0 19 21 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
317 0 0
2
43759 0
0
14 Logic Display~
6 712 150 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
43759 0
0
14 Logic Display~
6 739 149 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
43759 0
0
14 Logic Display~
6 762 149 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
43759 0
0
14 Logic Display~
6 786 152 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
43759 0
0
6 74LS83
105 650 177 0 14 29
0 6 5 4 3 19 21 20 25 2
18 17 16 15 27
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
6369 0 0
2
43759 0
0
6 74LS83
105 360 175 0 14 29
0 2 2 2 2 7 8 9 10 28
19 21 20 25 24
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
9172 0 0
2
43759 0
0
32
9 1 2 0 0 8320 0 24 16 0 0 3
618 222
591 222
591 319
1 4 3 0 0 12416 0 5 24 0 0 7
134 235
142 235
142 80
575 80
575 171
618 171
618 168
3 1 4 0 0 12416 0 24 6 0 0 6
618 159
579 159
579 16
147 16
147 202
132 202
1 2 5 0 0 12416 0 7 24 0 0 6
133 172
283 172
283 28
583 28
583 150
618 150
1 1 6 0 0 12416 0 24 8 0 0 8
618 141
586 141
586 54
363 54
363 46
276 46
276 139
131 139
2 5 7 0 0 12416 0 12 25 0 0 4
286 204
295 204
295 175
328 175
2 6 8 0 0 8320 0 11 25 0 0 4
285 230
301 230
301 184
328 184
2 7 9 0 0 8320 0 9 25 0 0 4
285 255
305 255
305 193
328 193
2 8 10 0 0 8320 0 10 25 0 0 4
284 281
309 281
309 202
328 202
1 1 11 0 0 12416 0 4 12 0 0 4
132 265
153 265
153 204
250 204
1 1 12 0 0 12416 0 1 11 0 0 4
134 298
167 298
167 230
249 230
1 1 13 0 0 8320 0 2 9 0 0 4
133 328
185 328
185 255
249 255
1 1 14 0 0 8320 0 3 10 0 0 4
135 361
202 361
202 281
248 281
1 0 2 0 0 128 0 14 0 0 17 4
323 66
323 65
323 65
323 139
0 4 2 0 0 0 0 0 25 16 0 3
323 157
323 166
328 166
0 3 2 0 0 0 0 0 25 17 0 3
323 146
323 157
328 157
1 2 2 0 0 0 0 25 25 0 0 4
328 139
323 139
323 148
328 148
1 13 15 0 0 8320 0 23 24 0 0 3
786 170
786 195
682 195
12 1 16 0 0 4224 0 24 22 0 0 3
682 186
762 186
762 167
11 1 17 0 0 4224 0 24 21 0 0 3
682 177
739 177
739 167
10 1 18 0 0 4224 0 24 20 0 0 2
682 168
712 168
2 0 19 0 0 8192 0 18 0 0 29 3
430 327
399 327
399 166
0 1 20 0 0 4096 0 0 18 31 0 3
411 184
411 309
430 309
0 2 21 0 0 4096 0 0 19 30 0 3
421 175
421 273
428 273
1 0 19 0 0 0 0 19 0 0 29 2
428 255
428 166
3 3 22 0 0 4224 0 18 17 0 0 4
475 318
496 318
496 302
516 302
3 2 23 0 0 8320 0 19 17 0 0 3
473 264
473 293
517 293
14 1 24 0 0 4224 0 25 17 0 0 4
392 220
491 220
491 284
516 284
5 10 19 0 0 12416 0 24 25 0 0 4
618 177
579 177
579 166
392 166
11 6 21 0 0 4224 0 25 24 0 0 4
392 175
568 175
568 186
618 186
7 12 20 0 0 12416 0 24 25 0 0 4
618 195
553 195
553 184
392 184
13 8 25 0 0 4224 0 25 24 0 0 4
392 193
541 193
541 204
618 204
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
