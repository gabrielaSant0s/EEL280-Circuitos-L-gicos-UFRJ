CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.499203 0.500000
770 80 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 119 288 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3965 0 0
2
43788.1 0
0
14 Logic Display~
6 787 450 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8239 0 0
2
43788.1 0
0
14 Logic Display~
6 683 177 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
828 0 0
2
43788.1 0
0
14 Logic Display~
6 539 159 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6187 0 0
2
43788.1 0
0
5 4027~
219 601 229 0 7 32
0 17 13 5 13 3 18 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 8 0
1 U
7107 0 0
2
43788.1 0
0
5 4027~
219 448 220 0 7 32
0 19 13 7 13 3 5 11
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U7B
23 -96 44 -88
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 7 0
1 U
6433 0 0
2
43788.1 0
0
5 4027~
219 304 211 0 7 32
0 20 13 6 13 3 7 9
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U7A
18 -84 39 -76
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
8559 0 0
2
43788.1 0
0
9 3-In AND~
219 647 492 0 4 22
0 4 5 7 3
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 6 0
1 U
3674 0 0
2
43788.1 0
0
7 Ground~
168 1075 226 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5697 0 0
2
43788.1 0
0
12 Hex Display~
7 1102 157 0 18 19
10 8 12 11 2 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3805 0 0
2
43788.1 0
0
14 Logic Display~
6 360 157 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5219 0 0
2
43788.1 0
0
8 2-In OR~
219 699 299 0 3 22
0 9 16 12
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3795 0 0
2
43788.1 5
0
9 2-In AND~
219 640 324 0 3 22
0 5 10 16
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3637 0 0
2
43788.1 4
0
9 2-In AND~
219 644 388 0 3 22
0 11 10 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3226 0 0
2
43788.1 2
0
9 2-In AND~
219 645 430 0 3 22
0 9 10 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6966 0 0
2
43788.1 1
0
8 2-In OR~
219 699 403 0 3 22
0 15 14 8
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9796 0 0
2
43788.1 0
0
2 +V
167 246 40 0 1 3
0 13
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5952 0 0
2
43788 0
0
14 Logic Display~
6 227 139 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3649 0 0
2
43788 0
0
7 Pulser~
4 130 184 0 10 12
0 21 22 23 6 0 0 5 5 4
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3716 0 0
2
43788 0
0
35
1 0 3 0 0 4112 0 2 0 0 14 2
787 468
787 492
1 0 4 0 0 8192 0 3 0 0 15 3
683 195
683 220
646 220
1 0 5 0 0 4096 0 4 0 0 10 2
539 177
539 202
1 0 6 0 0 4096 0 18 0 0 9 2
227 157
227 184
4 1 2 0 0 4224 0 10 9 0 0 4
1093 181
1093 212
1075 212
1075 220
2 0 5 0 0 8320 0 8 0 0 7 3
623 492
517 492
517 315
1 0 5 0 0 0 0 13 0 0 10 3
616 315
516 315
516 202
3 0 7 0 0 8320 0 8 0 0 11 3
623 501
374 501
374 193
3 4 6 0 0 4224 0 7 19 0 0 2
280 184
160 184
3 6 5 0 0 0 0 5 6 0 0 2
577 202
478 202
3 6 7 0 0 128 0 6 7 0 0 2
424 193
334 193
0 5 3 0 0 4096 0 0 5 13 0 3
448 238
601 238
601 235
0 5 3 0 0 0 0 0 6 14 0 3
303 238
448 238
448 226
4 5 3 0 0 12416 0 8 7 0 0 7
668 492
922 492
922 534
98 534
98 238
304 238
304 217
1 7 4 0 0 8320 0 8 5 0 0 6
623 483
570 483
570 253
646 253
646 193
625 193
3 1 8 0 0 4224 0 16 10 0 0 3
732 403
1111 403
1111 181
1 0 9 0 0 4096 0 15 0 0 22 3
621 421
342 421
342 290
2 0 10 0 0 4224 0 15 0 0 20 3
621 439
120 439
120 397
1 0 11 0 0 4096 0 14 0 0 24 3
620 379
486 379
486 267
2 0 10 0 0 0 0 14 0 0 23 3
620 397
119 397
119 333
3 2 12 0 0 4224 0 12 10 0 0 3
732 299
1105 299
1105 181
1 0 9 0 0 4224 0 12 0 0 29 3
686 290
342 290
342 175
2 1 10 0 0 0 0 13 1 0 0 3
616 333
119 333
119 300
3 7 11 0 0 8320 0 10 6 0 0 5
1099 181
1099 267
485 267
485 184
472 184
4 0 13 0 0 8192 0 5 0 0 26 3
577 211
560 211
560 193
2 0 13 0 0 8192 0 5 0 0 35 3
577 193
559 193
559 64
4 0 13 0 0 0 0 6 0 0 28 3
424 202
411 202
411 184
2 0 13 0 0 0 0 6 0 0 35 3
424 184
411 184
411 64
7 1 9 0 0 0 0 7 11 0 0 2
328 175
360 175
3 2 14 0 0 8320 0 15 16 0 0 4
666 430
678 430
678 412
686 412
3 1 15 0 0 4224 0 14 16 0 0 4
665 388
678 388
678 394
686 394
3 2 16 0 0 8320 0 13 12 0 0 4
661 324
672 324
672 308
686 308
4 0 13 0 0 0 0 7 0 0 34 3
280 193
266 193
266 175
2 0 13 0 0 0 0 7 0 0 35 3
280 175
265 175
265 64
1 0 13 0 0 8320 0 17 0 0 0 3
246 49
246 64
688 64
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
666 500 871 524
676 508 860 524
23 Resetando todos os ffps
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
736 374 773 398
746 382 762 398
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
741 271 778 295
751 279 767 295
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
900 237 937 261
910 245 926 261
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
33 21 206 45
43 29 195 45
19 Contador assincrono
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
